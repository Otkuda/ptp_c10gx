// myRAM.v

// Generated using ACDS version 24.3 212

`timescale 1 ps / 1 ps
module myRAM (
		input  wire [31:0] data,    //    data.datain,      Data input of the memory.The data port is required for all RAM operation modes:SINGLE_PORT,DUAL_PORT,BIDIR_DUAL_PORT,QUAD_PORT
		output wire [31:0] q,       //       q.dataout,     Data output from the memory
		input  wire [7:0]  address, // address.address,     Address input of the memory
		input  wire        wren,    //    wren.wren,        Write enable input for address port. The wren signal is required for all RAM operation modes:SINGLE_PORT,DUAL_PORT,BIDIR_DUAL_PORT,QUAD_PORT
		input  wire        clock,   //   clock.clk,         Memory clock,refer to user guide for specific details
		input  wire [3:0]  byteena  // byteena.byte_enable, Byte enable input to mask the data port so that only specific bytes, nibbles, or bits of data are written. It is supported in Intel Agilex devices when you set the ram_block_type parameter to MLAB.
	);

	myRAM_ram_1port_2011_wsr2yiq ram_1port_0 (
		.data    (data),    //   input,  width = 32,    data.datain
		.q       (q),       //  output,  width = 32,       q.dataout
		.address (address), //   input,   width = 8, address.address
		.wren    (wren),    //   input,   width = 1,    wren.wren
		.clock   (clock),   //   input,   width = 1,   clock.clk
		.byteena (byteena)  //   input,   width = 4, byteena.byte_enable
	);

endmodule

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
sdgfHulCficeOLG6pwBYndMfaS2Eo/Uap9JTo14s/yPgu9EPMM349dX+g5gsEQa8
aC1Kw/xnY+U9uHDyqzlW5owivPJ7kh/1B5bYlCPVroeMWXKIeHzdaE95uPphPXfk
4/z+dAVGV6l0l2O7AKXUXYCm+TwMvXvUPNGLMF64JpI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 21520), data_block
QJT3kEnfjLhk1NZMSXT1f1ozha8TSOQf4blX7u6Wajo9kp1O3clL9l0MK4xMq+kZ
pVLRLtd/vKjT4+jjogXUUSQYms4LiCuHrKd6LMmN7jopb3vlymqmBC51sll5vsfh
qUWiE4jKHwaHjJfWmn0R9j4Sjlo7KCssc6a9OId+UJKmuIcepGIs6x6RHn9PVWJp
FHvVGuxzgo7ZXxcB10MnYto+jZwETC9yG5ItATBu+j8CodAr5AXpRgEhWPiL+2a1
FlsID4+EeUE3blsSXa6Sa3uYsKbdqdxVXR2RGhfaBHy7RzmW6yDtaFs84az8chzi
ijC8+mi8Gcr7cxmWrizYWWxjJ6xCcyhLi4Ze+ZSs+67whJDV6T70tE8rX2B2RZv5
fZpZmgCZbGuVzYxO6iKus3vzyg1xD00fGISvGPSJptbyDoyLpLvFhf6XISt0SeCH
i4QQ99f+Zg0JslIdBd0zefGltwRE9PWpuSsPgCG/9uZKo6XmRhHLis0cQh0PBoek
FhxePXy/6yy6PVj5OWvqNVXddVrYGMK67zdIAAv2x8Zs1nBkzD+zTdjpEoZrbH/Q
A+vlruxkAOG4yJWGkzffs13H9XHEBRiWP6DfkZuEcPISjDWUCvWeswcPtaWB7/58
DZRe7vS3v/4ZO21b4h8KL/NNJXdA1RhkftJwN5fh9ahzN/UHT6GfUcAtNOCIJA4w
kV8K3SYOg6Txt64uNmmrHocxyRxvA08/ekFwmkw7UjGeeRHB9VyPQGgxrSPaoNLi
4yP988v7ZrlG4wbu5rE89Thh6QGACU1kc8dmUHaApjzZtlcjnWhTHu7lFBIdHUDP
y09e+fShi6a9yGWpRtof3dllxkgnm+du9FRPS3VD7NH9Zw8hHC7qdvSVtBgvpQlv
OwClCkwbVy5vR2rB/t0EoZ05qkxedqNNfMfpz6OxlhCiNVr7LPMX540LjKlfGv7x
Jx76eNV+NHc6qc9RtnVWlJNGq76R4c/LcaqXfez597IIJx8vXwbSP9mpGWNOvX5g
gqPL3i/sUBKSy7QborhXo/9pp5n+8O07LdKs7iyI8FEQnb9Qkf0kPpNtVRxW4XXy
WOEKjtNhCx+gyH/7MWqIRsWZnsed+4msk/r45jd/M0rAUXpqHHVHfrxKoYMacJH7
IGeJIpTNOSRWLdfgcXy5zFn3u7+ImeyjaZx9k8S4j3dW3aGA0bKwZe4a4fb/VlHB
JSpyUcZSBt/wK+8P7nTpMFxoVLvIXqCN+0cuQ4f6ZryG5LII3bpOyNQBk43JdB0v
anh6oUYNmPnW5y5qmxMVwVIHJFhUwa5gc5eoZGR0z4qvNHZuaSGaeq/q9n1UABjX
3IGm3igZcGHpgvlSNgaSrLEYxNSTVHLMrTX+2oChc6V1mMp3xJPcpHbGoxp5MgRZ
zsEyGCeGYE6rAmpreMMTDy+HrGCBlhtpjiAu549Ktfb4a7okGSqFBU1rS5Mj9D6o
HdF5GYH2kPo95MT0MDBJxP9Z/ZQi1bCWouq6ZD7WphxMaeY3RuAEhKOeodq07HzD
IxWFejFfZRYZKmbecqQs01FR6e0HX6tCBQnkfQqcu0ha7DL0QR/T3Azpt1KTnvyE
wvOqCG1WkBmGkT+Jzd3WKeoBhxBFMYcDTnThEvvnKcgyeU9yEskK9cM5jaWnFBYL
aM4ySQMy2ctn1J5Zb+B7bAXhrolC5J3yDR0dGk506xcrLKOJ6ZOYVq1NcOhyVo3I
58o/+6r0ds4Onp6F37Aeqz/hDomv/EB0gTPwcWdS+EewCDgvYl8zBupCaM5WFV31
bxOrRqoLtYAF/mfbO/iRUFTBlsKEsSRu1YpwGUIcZA7nhfAzLfx8bBWX8KXWcV6v
Di7o4jUjm8iBrqJiy10FV970hTgqMMnjQGGHbeXiHmGDWPsusugKggfhu0K1ZyDK
PArh2wkclxJF9DELryADiFrKyrykhhrGT1l4A8vuWwOb0/Xlm9UHFRUO6CehyiET
oimFldTOPTM2WUuN0yJqRd4YZOljvVcZiDXsbucXzB3QlMNzboukmQYC8PvZp1DL
KZoMsQX3dV7exrtLOiwl//KTlKkV7fw8ySvDZJYGREEiWmdUHbJWIh5eg6gHHRdh
7vNkjHZ1xhUdufbo+p5M2aBxReJExbp/0GWzeLQUd9lJfyCN5moBz7cXoernaoyN
OYNt/TY3Kj5oH/Mp7RHSBh7vXMx7yd7fKDu5zzpvbSSYl9FXhi/b6nhh0cDj8XQd
wy2apuVe35aXI0fQ+PDCNHPbFGNO6s+iLDWIXsW4inw6Z7GgGUVR6la9GGv9Gb1M
YKq623E+pQPV/K+6eJzHLWOwJkm+qvcLDYw1tHjYMbhmFo4ShC/XZpu3FNc/LdaU
ZCmPAZaWwj7es3R2DUwod0q9i5Zu4EoOUaI3aq7LFXxqHsc64MwZnDje8tvYyalU
rv7Nr8owj9pzJwI5CX2JxaoEDtdunpveYeEzavBZ9mFhTG5gseVppeng15JXRucF
JpYL+Zh3ekRgYRpPbaFGWIbDlOR/ChEJUkkhZWBZONEjhZPkLgkRPD5tr/L9niw1
nW3ldY2RYrB6Oc9IuADm3PYeDkpRx5DQPLjru2TeYNFz5rfSWOJr1u8OByrszmtG
ejPqqxHS4i7rpJNw36v9Gf74Maoe0TLwYRzH6mTmU7XWyrgiyjkbDC2Q00YQq3W8
oGPf+J7jcgPQnGo7orG09jJzy6UYD43FgKBIJsXuCZA4iLqdgPVl5W+dD2NEiirz
q0AN1IbAxfI2QOM2gML6av8wBJmrHBECfbbL7SBd2Bv1qFTUL4qOcV0wWnm9y1Jx
880s7I6kP0YLj/7MAaB14ZXHS1FDhQcbdLM/1zIBiy2vW5137w3asIVGtY9EYe83
bizqPz5W48FK42C1VN9mes874vJCq/ebe9Y37CI5Zc0T0fqBbRXK34knaFLo/Zlz
2bfOVdB92/XiZbTr8fLPdJFKTwaNjs4zz9oe3KtfvAR80HcR4lZAXHH3ocWkTV98
FOFWBYxQApojituEozhFnq+2/vB1l+lEoJ7CwRwNdZu8coz8zkyafJwG8/1+4f6K
tZRvOL+vskG9ksEweUPQbDtDwfs8Nvz1zriGixnLgrPmzNGtF9rdjpRJq6ur8Zjc
mOqkk2Kk6ZP/W4xn9nk9J38H7wlBp0xOL9plg3+sy0Ozjj1CQDKsUtBq9ZBgADiB
R/GXFmGE0OrkqfLidXFh9TVUOY55UIhO4MPiZZZOb49izxafL05TFGEsNQcCuwXO
XLa/z+XgVaQViNzMel6yB9RQTk0y7yCpbK1hZjY8bVR8saJfGsvC0kW576YUTXxU
heHRY1pxonfq1R2NxktQEiT/SLJtoCZK0N4n0Ab1C1OlLzeq1O+W8njyQGZL+bix
gv22rfiuUDlHggQGDvNw41ZS00JaotNTbDm/gMjfyTP9L1dxo+HOFLlqgcr1VZ4y
ADAXSf/HkHEt9YZPEOEmhPBlkZMI/rZ6k7iBEDBoeIRHqNgsmUoKEX37W6PzJNg3
dK7T3WuLwtB8v1kAOCLpt4lUFCohE0WYNYRbLnapUrrnSFBYQvfotO8/mFfB7Oq9
b3wIg1tHslSJiCLPonY6cKQ/GKPVLPeddNYLBZe3sLzFTH+X8HYv6S8crvlvLkJ8
+hB/5ApYgq+ytpr5nqWln/QHLXQIhcpJ+7GS6k0K1ug21WvCWlhj/BR2Yc1fgFzP
TL4iS7aQgrPzDjDtKvNd8UZGcHNfCvZoCOrCLu1XA7Psf57Dfd3te8ZoN/5SvoYY
LDKwbR3m5Qr9U1HWa9UEru9YPwQYLfJMgK/sTICrOxJihlp4tgavGEzk0n/tdvs5
5lrQF2QVDA+1aXVOsJxFrgO1lmbywmTNp8llvYxU+zz3q5MUP5ev+GHDuRy5lyO9
pvLbNam6kKbUcxIPxDWkjWEKOw2OKNgkrGP73lQQ81/m0scWWHYDpLoHh39woRmE
zXwHuodXmGn1uqDPn6CCEl74/oLnwKCrLpYQ11LFy+/z1jQQfJaQ99Eg7fW0zjnf
ctvuCN1N1FGtTivA1XNtigzAzPOGabLiQN3OvQD5pnSu03dKZE/ICQvevdNBkZPs
RI7ZK+DF99YkG34hvB5QOxb3TnV6DyakDoaTi4b0zAHpTYKrJrr8kUeBWiNdpUAH
Nt4yryYihxVZE009UYLSnrO9tSbQcc4npob4T5MsxQzTw5yK29vETaDpJ+FXWHQ0
URCofXhhyEvvzBVuYk7quXI41VEi1bf/9+KjgvEeItma3nfh49Byy1JQ2oyl6tuu
mH5Ew0V/H4CwfjiktGW9hz395uGT6YUCslgQgNPMhZEJ8JJxm+ccmo6XlJRXbOzl
j76/xrvNMTD68FmoAAXnNpY737XBrxFeDycaaIYYI/u94qBbb4eQo6GHfA19MbtM
ozWChPoRlzwd2U4CZLeV5Qi2hkZ64rgEGV/3Nug0/CSp+eNyQEjevlzqyYFn5LrR
3YIk6r71MHDyg2UcBDOFsZXNuJK7HMMlKdu1UvCOUhtP3E1kjXmnOLFedMRVsHpS
+pOENLwx6s3kPcXH+7HLsZrHAdraHs11Q0UB/B/5jc5dfPiCzUTzY3+hQd5pJDk1
iWETHUHrIo9hoPGjW6S0h03C/yMj3hLtU9oZ6/ywRyzf5gr7HBqOp5KKX4kN7EOI
zv3brXt/TB//hQWi8N1YCc4WkddKXkESzlAqK/F4SjaHvGkc7XdF0To88xnmIxdH
sr32uAVLQg2Zz4uYL/3jYfAr5x7HC8xzEQ8cnr4Ag9BgasXiebGIwprKvudnVOK+
1Ll300mqRW/juGq3AuREuYuUA7YVvRhUM8zzdoQvkYINk12Az1m9fbvDAAjsCKhl
XA3PDWDjy+EbV7WFgKtTtK5NQIqrhIYJ/MlNpID5pmPg6VbtyZoa8iBTVDwaWcll
D+YCWpNmsVXwx2tNsOS19If8uGP99I8dw2eulk52OjjdK4t+71YDDgSIxlfGjAmA
+gsyomLHh+EhzL3rxlmYpVM3S6Ti2CeRoS2VB8qtLRsGUyG42oqLk+gmEho9PSR5
2g/u5+uxjX9vkEfKEuHjHc1oDbAmhhYIqPNgS9JjhfYsDIuyzVZRih3aKzze4Xlp
uynu3ELVrghyhh9PixWKZskJ0zGv+TQrauZv7T36z7B0mR2ZEup68z5WI7hyI1tU
3jgQ19SrTGgfVIjdRCIvcj6eICXKzt79s0hIyRcw2vZUsEHPSyK6mh/s6CHcZFBj
Do01AHXl8lZjv+F3XcrWEG0Snd+qfxx92qIceeroEvmc1WEuWka1rwOGDw+Z/6Fg
7TgXfnpp/tOgyjck0/xbK3kqTFmvW5HHWDwrWLyNgzkK9NvyevYj6Twf4U95yEus
z2p3vGXCYdfYaQP1LoPhfUPEphEscxrufwWwzV/7CfDk4iB6t9042ao2TWR/nwnW
qLLHZAWqjgGFaMFXrW+tb8oApkVNuAbT/rLS51NWYsx7qDYOrmaNMVgcEKiLQqLd
CtHSgMUWyCiiW7ZH+02gd66qUZ7jViWpcYxAUrL4u7rABSRurFUMqD1IKZOheFJx
p+vScgYakzHMETaZBWml0hJKxz5nPNji3LFlqtYl16fjTOtGWnBZgCw4gWDcov6B
Tg/I3x3xrx1loUna86VFGjGZUBVvegkt8THR962fC57/vsksb3MWfFSWB6/l+0ea
UX6KmEuOcPRY/XmgyFgex/37HKMeQnW1xE7oGQ47ejnXom22TGXA7VBOdv/wg5Qv
ja+VUWxOD1sTQ2ua5Ew7LMyRkNy3hVAiNpnrodR2nULue4eZl2uJiiLRNrRVN6pr
aH1SVjxsM0XP5+VMX8JgbH+L8dCOiUO3wIeN9ZGUrdEkPui009CmqfUIPHLOqJHh
VxKAsphWo0GWUk5zEnJdDCo8bykOZzbChCwuWcaA1D5rGan00u4vwbgU3SVLY2dE
jGwnpm8Ry/8HZrH+EQi8zhPbyagslQaDDGxDgJ1/wAWKyYPHnjKw+CGM7/OA1G9D
CsroilnGyPjJN3/3XQ0ukse9kBAuOx3smsrvG/OwEls9MArfdN3NOYJC9iU76j5L
2tCXcjqhKST7wJXn5j7d0I7G7nF+I2zaqOAZMZk4FR0BCPRshQxy3hACS/J38peN
Q9BDsXQC6FfQCwix5bRSGRvIHm4O6mr2L8Kx+FtsA4zqB/HZhDHUQarjyZxnI+Tv
E4B3CHJSQxFR3HXn0m7UWrpmYKu4TzSReBfK0DR75H20qnkP8ZHRlTiOLSfodApM
7Sz6Z2SrKDfceutz6XHlVIWeQkcNfnzgMlavAqo+3v6X0YyKFJvoETpVKT+1pMZv
VgceTM1DKnqkV1ZEAx6TYc+TI2HAgCkbCx5p/D2ZbenRmYuLmtO+9IWW6lyNpH5Y
8xHFXZUz8mmJQxvd1lASPVjoIsdGiIk38977RZQrQDL42aDqboYNliIqjd6jF5DD
IdAem/LoUP5+HyLY7l9azOpVw6SkoswBRBQCMktl6oGIJJWMH5xrUcUG8g1z0G+B
wzKKuMvIH08hMGZhd9TSP34jpeiwTSqZhAOLAUqsP3c3p0d2S+qwSYYc/ESJuhH2
e2+LGXgro99bGED3zObnWezkMvem8kqeweKwz8lpoiAMboojTSN480PRYkoBQYJU
bdxn2Wl60plRBwBJ5ysDB2scroczTxvd1dB/06buNv+tSPB/SMpLcFvaFqJtdiYl
6ewy6AvtiJapmMSR8B72fOIjmdQb5ehEuJwg3OTZoRZZE5T6FVsI306VUHGCnsHi
8uBoBMxEjOfrmxx4Qj/B7VXpNcl8TMU8B8Owv6LFnUct5rR0uBSAErNuGWo+ONnx
/Z3DxxejnEu05WclEWYko7two8VLEnVPvP8lAuOCjM4Al+OHWYfdtRaf8Ym8ROjR
aBr+FMR7BVvatyJEgWNFX4QUPKCo5StxEiga4hkOtFSxlS9hUm3/jnWgvvLCX8Si
gfPntEj7i8DPelGcX3GAyz1P16wIpahr7RpxKUdBOdgqNxbjqcahQ/RyDbzYe6X2
zg9RX8O9/TMJYUD4FBEGoO8nz7HdNxrDPsc7rDy/tmNtn1xwJ3dgA69To48dA08m
zIkmuC3IHzhHCPyz2stUfWFtrK0bFiPLcLQrjkxn7ei204YJxewsebsnzQtdNgWD
b6VVDpVzWDs1TgbEsYYSFJQ7DrsO50yDfzTlDVoUggpTJeySxfiR9gKphnM0EK7P
cZ16YGhRfqzsH2KOOXsECePEWjiz29yZOJJ880+UimbbWPxPygdc4HF3PEvmdzxC
TxZc7vRKLW7uulszSl/m9a/GIedzuLySUEzY6FupxR9e4+ZYPcsCC08Cr/aQZc+Z
Ije1CF753tsKt4UMKOc9C3Njl/VtXo8bk2RnTyj5cmRRUemKfU1lyIcV2tTkf8sa
p9xWM21uHc+Ra3EfqD0pv0AsV1oI6O2n2Dz0OReN8X8fSb4JOfE5jXDHjPoXB4Xs
thcX2szALZhYui4fEVoWv9WJ36U/sTc5UbV80am4lHxRNm4whUWMextViHafbp3d
JA1yCzt1LOmsgDLSeFFYbYnVrcn+YuqknUFKXlqxtfGScADH1TGfDWnmfPg4SJQD
F7NzaTaYvTwGKldL4BxzAlAhsmUSK9t2S8aDip/iEIm5X+N4g3xfHffK7qAiRBlK
6kIR7ahib+EC3CdCOnK6VAP9QrqGCpLGzsKp2Xn9aTjrR7EWODkutuU58WD6jNpC
469L136Q0QEl5/V9RQNhFQLvZ1390Qz0QCTAbK/U6d5wN/VFbO4mCcTLvPCEhjCI
OPYJchQSmO0enyZ9Lw0pEuKRXI04J1PXzfYFU76LALTp8aZ3w2nJ5aPHkOXtDyUt
H0YLJk8Zg4eWpTMduQfxf/fDEqVXVnhSGm8mq+DwtR17u7Ha4OGVeWrLO5B6RSlK
NqeDLfeAMdc2ONSSG6M7HbMPRpopEBW2S/I3dPU6UyR1w/xKr+pbEW1oZvqMA6PI
WI5UgoILyBn/MgtJCOwlKUhhdb9pKAJL2rLk739LOQHL6SLwmG38Kn3ufWEilY+Y
hJf6kId4FIbA90U2SMUPAnfhT9tqwixrhp/rq5vGKwS/iZD+x1IjYfOL49MTA0fC
YtQGHHTeR6VChbve38EwRpcoczNX6P39lbNtcEoCYNt0vp7gwqAgf2vifboDIDUP
AAAGJEnzllpmYGP7862B9RHzMz1PxxGyghrnoHjsVOCMLcaYICnNE/MzZU6C1zwf
825LYP/BAp82CfaoJx9H7xH/EA8c8DTWnVHRLTkC7cL8MH7Vhz0igycGg2hsBEq5
2fwmwkrKN/EOBWKggrZ9G9MYBLGzzp0YtFvyKpFcKo+HPxhQtkoMVbAO6yQUPgrY
PdzBYb62FGekDJ+9qX1Cg9b1FSXTO5eY0eOx1MPMMq0iGETucN6lEK77TW5bjEOw
+NtDiRRUCxIrUHD62Sns1WzXY3PH6wiBubg9ZpXX/36JtpTDRumImK30KNnjebju
2u3dOV3xgrAgsME+3Z9tnNUppEvKlVUUPDjmJ+2drzreyLZHwkiD0uRfLE9eiCra
3xGX0DDlrXgOPDZk9vPWtzE85J44dVAb8rcDFO7liJgICy9I95uDXBklRsEuN14A
ZQHXiPAfJetnyJveE4PM6FzqQwPJG7FXZIKGJtkAwkwyNF+H3gYaqI//hyBswrMO
YMEV3gORHn0sgrnn3/5fGzuUXE4Hz5ITCl/bFZZipkn3SDcu2+4xdFhXbIlAgyju
gN3Qn0stmxvTtj+BaMjFSkpZr03H1OmDWi2BMRe15fBl/n+cp5VRf58fSS8zvRIT
nvF1Za/CN2/w+RhMPQ4yi/6EoUkMck3purdaMBTcUwnPVyePLoIS3L7EZeajUwvf
S6N95YUlFk73miRbatT1MEOfP/M+1Qf5lc39QRW103P+/PiWaFWQrw6e5bC3kKmM
F7E5FD6onLzQ4f3J3XtDKla2FWNZvYNbYbzlJ/rP7tgOg1IxPl+KLJjqIA3njsbC
DvwkPh32eTN/LrnaBPQVcZpAZMjioCGKzunk4O9GhoPG1JTJvu8HitfFPbi1X1DE
L86xCn9BFu6cOVmCGgPDEcXSIejmbjlPdGtRGuH0fgF1p99zn9HSK2t2LsK5oCND
7KeUbVFcEYFPQ/laATwNjMgzHY24HU75yGs7fMZ/QaP3MvWK++OFTwcXuFJP3Oym
ew9CcyyQ75qyMRLGNwdcHLfIsm8vtWa76qKFgPJFw/n8Ruj8piQhTsSDGBj27EAI
t1tfqlQMGMHupbE5uCOP/DH7gRNbGCOq7m5X+ywFWWSxgS48iIoZA4HrP7tsXG+l
/coheGMnq9ZTYgz22nHyOF/gdbVzottZC0J9TPjeShnPr7A5dpyK4w+4K4Qbb6kG
GfBuMpwEFnugawrxWyXV/e5JedrQ30pLMnTAH7CL8h3LMu1t3vSjJFrJi95Ou9mb
50iHGt+7/PKAmLBUXVK/tya6MOf/Iqay/+JNQQVexsbKmBBJYfRCo6wOfeBuc35j
EDCWRPIcUOcLbfgHspqCocl8BIevh4p4nPcgOmWLVBZWRcHe5PJtPXT5gsUYzlPH
c4vBdvNb+TmMimDQSZ0LyRf3wz+W8m5ucnS640HItfQT8fVij9nYKpzbxjsyy6RQ
24NvIqjfVxD60UT2XYzxIFZmaAjhe9XJ5NsRVDjFHOtA71KvLyvONqBoXKMll065
5vIykbWhsHMrakTWv2Yak9XRn5L87sHzeHjXJFrJqO6BpXpE2YkSbytukHoEiseg
pudX6SAnOeMK0jLiJ3nh/i5y2bPDcU4/8s7aa/8/YBvXKiByufTDNprS1fZIEUpJ
aYwcEKueDr3JrmPV5r+817zv9g+NNzu9V3a3AzgRePRJ8sqycTg9xQHvIrgAcp4F
JE4VloIo9t/8fogIPuPYogYRlVqA7QJhV1zwNEXLtwd0Hgj7q1nGf+2FhdPJnIar
2/bLt1lkleVLrk2e2nFzxjmNh4I44so8pltES4U0pA7f8riJeyzbxvFsMjpW57Bb
wILWxXMRP4JlR0ieqFpO6DUvpI5zfYeJ+U01BzNUTn6RR9m3TDBFOy+49Y8XMT04
Knyiw7ykPPpH+aA20XSEo8Tup2LkKhE4bUFbxghS3Us8VnoQFSuRfhaaZgTbWQe9
9CCGwyz91sXvC1rU63s0sA6laYxmFGy+8cdMkyvS1gXYBpJphp3o370oY+l7Ofvo
4FRbkRGTikpOycbsKTiIR7MsuZsHuuDGLWgsDkzo9OqeL+XsO4v6+HHTvxSJHEpS
l174WPwfUNpNoDrsO/HYSosy4pkhsRYpfQKzKvHj+BECQfWiaoC13n5jyTMWYKQx
7Fkhe2Xe3p4kyCmQxbpRB6wF9NEEOH7DfVk19g2/tdbP+gWC3ffzdvovk1LBBW0d
7ZrGxTO/xla8rrA5dJraeOsTHxyRam1AmZ2Jt6jkwX7/k1JfD9T3XXqujyLoTV81
9EOzrUrAn5xZMwpV1iP97SfhIRiWM6f2+euyC/81cYwI2XkQFgDv6KDClh6dTwD/
JYm3HFGdfx/yVIBNjLwzJfpLRQk+uPdFh92wUrdu1cfpeFTDe7BiVYWZQ4WpfpFR
rbOpEOfiltdKqfIqRF+PzKp64AdsXB32Irogr6nzggz2jfiRBfoxBMRiidHFcTKj
VVMsfDHYLT3Md/hGy0IkipB4SBiMrXfsJbkCVtSg3J+Q1BUeBQcaBnTVeGvibrY/
eVLCV9xR5ruBJU6mVSXu8RkZLlDvvX3f/PJDnDKv+4ouNvysP4rNox7vohUi5auY
OVZao3+LyskQgZJjHZKfRJ6KheVkGiAUs4GbhPaQYnua/VXMsi/0oPm8cdOVD4Rt
b02dSzSNXQ0YUfCfdWXi03etnEp0c9CpCFBVyFtPbtrsyGdi1Wo8IeGk2NLEjYt7
yNrD7NDHmOlM6RyV2XqCbY4eTB1V4XkYEWOfVfGhprtDDbU0gme5lmNn+nba+yF4
wd7afqJQaA3A60/xVZVpzrcF9T+CxxPPMNdXoTfUsH4QVx8r6hBFOJGJSru1yZRO
ejhqEeWIagIlzpraPEmxWIZmAeQYcWC2CFQHZtLlpbus5Of1+L5HP+eSN8DhQ/CU
rNf0PouHafYiWXG2IUdhyIR8msFXbvrwyYlRb/F9m/JTTwnFVMspHm1okEPNV4UV
fa+1vQOjBfzdcy1DmpZTPZLdBNy1LhILreaC/trcSwl+CTz8K/Fmc7TShG3ycTQw
Yh9a8ITl7j188ngB9mwBzDoKN9dTUuveV5n1Ud65tMfb2Ezx1AIWlWuWSKIKG9t7
M4LmdN65bE+5oq7LLNvwd4Q3bXYEzZqYlCnqu8oJk4OFq4pjKqfgZq1ImjktBYRs
s1y0TZl0KAVgN2cQNXil+6n545QbF4gLxH4CU5FrTd7R7kdTmAbi87bMjszJfB3c
fNY4V7PNjq/Z7PG7MqZhjytHr9tbfQ+MGzmpSBDLsyPGde+StslNgIqnVDbY5z3P
yodgBR0nPFYNnr6Ha5cSA+ZgeCJ6FYpbtkmXaBqznazdWCWsYTinhxspMzZ8v4dg
SUhEUdqXzrmxIhKUT8re01NYs6PslsKTTZ8StNaofpMj3AQFnngDrdij13VHslEK
6uk1DA9QihocIvxjrlDZoaA5MUVYoZbcBwwMlZ3pDnHrm1tQ4vOL6FhDZgcL6kKU
u76OCSVIfDLnwCVM9rjwhbiSLlG204rqayf++KW1Jk1oWyHzhGeqoWB3musozGu0
b5mWSzd8hzTlWIzQPB4WV9jLoNd7vVhyC/yl9dFINM8OLZmJXDypCdRfS+mUgH5S
ESaxBrpA9Ql8wKbiHyVhleJccApYJcjgk/85jSRT/AYpbtCu4XJjZsF+HrrWBlgs
4ICzxZYIntIhXoaowpJvkPbUwEFKc8YOGqac7b1bDHjynRrD3jALn/CGjz7LczrA
ILUkbcBsAvGp+zGdxrmNXgcypD8kEhoSmWwZBTIlg8WdzTJJ0mIW4uj28WXhr9zC
wASpU5xuJZiVUAkmk3J0wtkrxl8hhypciSCc49rwFf5JkNZetObyx0UBMX6V6ery
X8NVS0w+vDhaV4qUsdDCjCOk+l3FDX9LWiGlzg0PZ64Jq2xHZ2EVARkAFqounsQU
Dk8t2uJ3VjoCYTrx50pTUXJpo93WlcwRdlw/K7YX8zLn2BODeyMgKrjVZNUBaL+k
7e+0XqsRW6AV6Es89tyFyUsNtzfY8aIIjEvLfI+CUMnPw7PocrC7skEYZfGJETQX
4NolNOrPcL2/S6mWHy2Ojs9OccaoMUJ5pqzOPXnzZcCB9nWIeVYiiPIw7gOWdhws
f4mFI5Xp19T1qgc9HZ9/Es7QnO/vX5W+K+K0HOSU0s/XswxXb1aleKxITqy7fCIP
RTz9QxW30SVPyJiuryNqE3MKevIk4SftbcA3zhcfZUsLVK+3V2MSYK5o5Tyt+kAD
NC3zGhUteMp5PDA083oT9E2yvQPzrhxg3J4kDSpMn7S/gbr4uoVCObQKeggcDax7
Tzwg4s5EQUySItYrdHQh5C0uuqbIXZYROV0AC3EOFLi44qNVz9vzBpSrCBUW8uy8
sHZS0lnbrS9Y9lxo3Pjhf47ZFWNvkjMXR/UCjGUwdyC+HDqHRXJRbZ6rXg5mrbOt
6Nx1szbQNt+xObiJ2r2S/bQbOY3tcVEG8tWyjBV1+HQDouy/FCu2FriqeC4EvwbJ
ec6PFiC0vIzdwWekJGUhLc0yo3nHM4blAlXzDiF5lqhJzpDosQ6c2ow1q8topboZ
wsJuqcRr2vDSz3Rv+aCqb4eYWteLKIP8ckdYMUAmszeJIokCip0r+WTWSjkCw0Rd
4jnB7AgviQR4KzQaSlpuoAIcuyC/4O3RNgxDFnYm7y4H9MRm2pgG7wRVDj2N4Zab
z0/eZEaRw83q7ol6KmnNMkdRl6M7CFbddsV9vxnmYlZz8fSyUT5kU8UFwNVObLKi
j0ypYo+lH7kUTiWJkvzu2q6XfpKVZaenze22HMeeYLkp6ftpgT2E3heaBpJfcuCx
i6Uy/MAgOjhCcni7Qee3/YMG6aFzi/ipDc/V9opAfy8AZWRjvVZKBOLZiCd8rH9e
k8/96EoDLlceVU6oW1NIwC9islblWOgM8P7+atRqsiQ6yRH4w5p66uHHgbP+8F/V
tlHy9d4RS7ZPjZBpkyK5ybZGej2t4nAf8KPkU6hdiNHwTa1lM1xjdtgpJyU1mOPv
pHaagfMC4EVsEqJWVg5fjII0r/h87skGGtHALYJxLtP4BVKxe7OqCiEGM87zvmNy
malW4e3iE2buP7Fk6Tk3LIQZyyRFSEjHMnTS/Yl4GWGHedszKBLAuAGDCwvorYR6
d4F+guriX8afnwfmO4TJu6zBLzF376igbJgsb64IoNXOAb3CH+afLXoGJThEHHBb
z+OxbAxA5WwZXCyq0JEIAloIIEMBAjTbWxl1Mbhf7LUIF15xcVoxsLwSSod/xT62
nROTNNztJ2n4HBFF0LIK2dqzUgvNTHkC7jhhw3rdX97szy3BEiyF5D8ycNfmlvyV
vN86D0gGV2A8AOH+fjfgHhjXpye2A3SAIREGBjdEMRINFGR3wUJ0KkbVp4puG0I/
wCBJlFSf8dJJ9UKbF4cv73nfrhJuccQcXCBA99NJf418h9ZRDeTb1g/UAQcIZ705
3K9jss6/vNrynD3HlHFfj9dariTFUrU1LCzyqm9i52wlAmfChG4N5LNyXkzBOTX9
2R6vwxSb8rf7K9iq7ERkVEW3D6FB11xDdxJkQZY1uaF/DKMFStBA3j0hqB5iawGq
VlyQuZnsWEj8mq5FWB0EUxSskPdV1+NNuWeWH21gWaOyrJskuHI5MUnjewb2ocYm
cLMvRl7MFAAeOvebjRzvL+26y6H/rYS4KpNcEFYAeqgZRkDDBO7fYWUetQt0qyeP
/ezvPM9IlKLnPbq9r7UTFCEMVh2ImM+/inyP7FLaN3rVjmOLxdOgG0VS6jbPz4IS
P9qVYpP48vNzn1n0AZdpVjuW52BKH1bSYw/z01Xa4gBsM90xvP4Xcr34g1aP8u1S
rWlt/nynYxyjqcM924y7I/fYCtKHVQ+vPNSq0j0sXvfWeirm+PxceKSiQNQo9RX+
PwLkCLwmV+J3OTfnCelEamjnOYBw8jLBA2JsWuom+EwgRXOjywFk1GEQYYIicXeL
4KBFTeyHyLPit5jgJHLnXWYx4Zrd1zozpVPEpUZDHNwp9G9kJbuZtqmdSQQEzToI
Ginq52uP4E3l8L7F6qi5i5zLaqWON0PPR3zP0PUr+OAVjumKDjeQBs7db/7zBvCv
3mRZfpObKniBvr5gBrQDfLmwXkc5IqMPUbPlHi7NEqpsimHmee/l4/EsDf3VB+L5
mtVgPtCTjWE1BQaEVMyeWQeAAVg5fOtiAV+vyqwFqeFBhEAvzOeNNiPLB4KKxt1/
ph6bzoJPlDw9JbCuGyno/lzbq2gC/AGJvrJq6jR9yx4J1GNuOzecZRU86+NdSQch
URCOVJS1yAdgYz3EqFGDUl69ObxnJz4vtAG7u9GFwW54IFAHFxisDqokbshlmHJy
mjMwo1+/32zZIklyh6h3hJUU9VL2cB+zEiusa2SVpFjj0x7swYi7HD9WnY7rdalI
Z+0ADXLAWDcWyUMmCG/wpqWRJ46asH8hWHf5MC5NdR67+eJCNBDB6SiN1AvVBD6R
2xEquU/OFcerL69rdNhWrkBV9ifcboeqDsZNWy9uJnvxnKNVrneKgfbjB/nNvJ12
KtpFCZBGDyJ1VXrtd4wn/D8sKxX6vANcS1W9F5ql1dAeB3avTMXezdAzbn0LtxLT
EHxx+9mEsaHCyWcmJUXy55tHEs0GktDajuZ4oWXAW4+YABMTQlq6sJUlaAYyqAy4
0hag4TKD6G3zzuEcos0Gqa7t8H//jteWpA1AeS6sfKu/BuygPeY6NPSwPBr8jlrc
QvvZxuRB735j6bC5eJ/Mj6gwU9MXneOmbjRvCxKIBtr8I7R3adOKtrCUb0Pi7yBd
r/VBryyWhamNNzfv1fuS866vdyp/gAiNfEQIyuvWeSUKO6CJ9yKfFeLUYbO6ed5s
TtNy3mmm7hdlGMv19E1fp28e/fGiYhEmD5bX1GNsGeiTRku7Fu2/gIl0asUFeeKi
XAk9D9xAmpPfxV25hvBWvCLBVTwMwCnpfVv5Bo3qvydtRvPa8+4EMWyV7piVmPbc
SIQAK3nx4k2u3mGkyagbNIZNnxpxGkWrxTjeCLCZkRTdo82aDvrCGXhLLQVkLfdR
Xx0zrjZdPgqq5BA+nhpFAviJrrfayeV9NlGUTOmNzOR2Y1ySemvyt8eMK3VCfNtK
faU0kUaGO3t22isUeGQpc+7CiIEnzAk4sFNv45tkY+1Z6oLnFnIhonbkRvyeJ5Ty
hBzA81enOfuUojp/QF13NzeOakndh6YK5YS0sYCNEYnPw3GgAlcOoVDBEcXynnTl
QNB49LkL4Uxp5PzA3797X/bJ/dEc0FZ4w+FygI2NwoyWlMsj/DN89l+erzSFW334
bWfEk68sav/x4+HRk8iNgbo9IJOK0498b4dvKRPJjaJFk8Obw5fIMBiuh5dpjgeb
OkecAf4pB7XoPcWxwADwegGqEtHYipzsn3UDn/Sog1ui9o4epVNYXQ6mvmx4KwwG
KG1qUruFSa6z4brWH2jVRWc1NhkkaAnZjUg/gBTtTsCZZ1Jl6rMkrabTcMB/btg4
dLnnuh1GT+HsWnWqzLOv5J/Wp0Lv6Fw6IA6LFM5w0N5Sbs8a+cVRFFSlD0DydNtC
3YTo0UFbD44nIlq5xqsCqHIRCoM78Awbx12aPAaHrwrC0ErPXMBrSrLL1rkV891d
R9OiNxkbMp755bpIT9ItxGR9lGlQRPvzU3K6BoFBPpG3Y8yOBtrnZLvXaOpSMu0N
9rJU8XFIGdeDDhsnBdhAq3ThFY3nK1kHvwoksHspM6SjGQjXHhrC/SV5EoC7kTGc
0eWzfDBRmYp4DPzjNxwSOaF1KVyLX5ulQ57a9ehC83NAmzRIHUJ2Xw4yxnVSXMTa
xQknulHBZZxNTJ368ZwO3GhNHT1wbfE4/jsj7E2Sc6Kt7IxjvsvkVcyqcPTe3b0u
b9wL23P36jbhRHYYNLgYlTaVXGDjqedauSFqNAYrNYm/+d5Tj1txWXaymw4EIL9h
9OaLicdsFGUJcZTIFwI2HyDzOlqkD2dZwMNWIAut6DCGgV3aYXpcvpoaOvPbbhRW
w+889jfQcGJch9vjzScjWS80zD2dAPdVesSHfJvOnAHXZ8mrr6z+l1OKMy+uEfr0
gN64qpcdyIbd0flhNLP6uv3V4cZw+XPLkhZfyW/7v5l4vrvVIQCCQH+DPgqNKxYf
kwYv9Y+IKLNsr1DnjMjso1bLmpayu6qNrzf+Cg9xE5jaoxzf5IvfODREkntIHxCJ
G66xEfDto02M2fNKBBWv9u9JbEl1V3cqgbkMKBf2kMujiWoijsLzn6T/9XRU04WJ
VKHI1ICpueYfmjghoo5x1BxjRnSBufHqlC+bGW/CcfnWVPvX/zEiPH8ip6XJKJTe
lBwnPjyKBoX0hnE2iUloOJOLRwhgXPGMS3cnbWJktKRxARVNQ6PHWYL7tOZwaVmP
Ao3w0tkASCOggNDFcAngMKPrBA0h4balHN64KnkG8p4yrHGnnowgIRfVSuIVfhSd
vy3IftrfLeY08fWrhw2QsRnWOhWkVEBKsKKc83vLUHW11581zd0B/y/gIZwo3fq3
CFZgusqAGHfrU47DgU7GvO2iFFSgpfA1xJnFuIN6cblx7XYEpHyzQK+6Oehs37dh
f8a5m4pXSx3zQp638WkD3xA2WDDCKWmOkTR8q+lZ8exVIuMzLmK3ny6Q3HCbdnTn
2lEB8JXVI6QaGgA+1KDZLToV+odiXqDb3Bhv/IQGTCVLZM32ryI/91xNBbD7Bmyi
tKMalXJCELHo553AI2SgrjNbMP/gtv9bwYJNLwkPO5uf5oJRzvR+Plsxnf0M1zv7
MNLyMvX6ScnrY1dQmrDzA4R+LaRRhdRK8+3P9eP+pWIhnvzEpUXEL/T1cfDoqEk/
IO8h+y2mpex1cmsEMvFYTHHIfk6bevmYjni7rxQr8u5UwX8MlkcOhrCno1Sc+8sC
lbE575xNnsaUX/Pp+QXmtw6k93tJAIeleq6rDXDwcXuLBIXFLlA+sqM3vKmwb+84
bUZSRLyBv+rLrxzFPq/0abSJk5G4zL/wIBGJFPwE7yWsZaE3gnZNOzx9h84pZbn3
jMq/t7ejh7Y7sbiOL8J1cSF8bpPVfigqYVhRE3e3Mj/WB1fRDD4lbLCrLcKcM1AI
2Fl+rm0ypupoe4dAACUQXDELytFNdeKEM2na3jgqSilq7biw0L4Cey8oii6qRD1g
ipJ+Fuc1PYmNATTxnlQ8oBTRnuCPLI0X/llwVIVDwalyi/W6eSHxsxbChzbAqC+S
K5UqFiknf5pXEd8AB/H408gjUWV7BFT40nLCF/tSJi7PqhmKCD5amFQBTZkbat/m
uvYN1zpNiMj8ECMKWgGgc6Y0qZxaU7WxXTolHlc33uRHOC636yH2ShAIzaaMyYAi
yNB68gH32LVmXQ94qvobMeV0VGOxdEwfHBTpIuL1HJfblGPPxqFR83cfh4KISKok
8Aga1Y9D6t+WZ4KbVneKvxqFvJrH60356kDFWm8JOTKPQp4kFfucPzZBuNJvR+vl
NntrQ5x1IS+Y02lGla9GJiD2loleO4BQiOObCJYArfzahDMVPMEl0j1Y+L8/itqP
YNTQ7C9svecBxaupgsbEoqHhAD75nyndPtEJwa5q4WcTJr25SB3yniLg5RRki8MF
nI5zSJWwTK2vAunWv22thvmXteHZqU6L9PX8AkMEBCbilEl5X1JnwI7LNwfgA9Fi
Lzj5NzNdnCx4ZVstNtPupmau76sGuhxCIQX1zzqtqxus4GLa+TDksbM4Ncwf3aOe
DBPYBCBgIItVHuG+n+L/jJjdsDknyhdfCC++hJWzDACF5ngf7/5Mdippv66j6Ej+
s6YjVjhgd5oOPiiHoGeSiQ7kl0yS7nzvNPiNmedpQwOJR2cEhz6Ih2Gs6PaCjdA+
9z9tYobL+WeEiYByDE4Em+oLc6YO88kom/IvFlcbxXBgXke3X4m6iAmxyV3IMhEL
xTZDYf7ES7i1XylZ70g9trMrC2iqoHXVISQoOMgK34ZfXC9FYRBYw6LxVOBSpAi/
Lmz6tTRnp9JUTHRDixcWTGuGJB5WvAfEEIEFji2fYGwunWlH+Ny+yUkGB5AH/rvI
NybFTsOMpyzZXHAbVvEvFYEHEdb2oMlBDb47Qr5ZzhGUMUropJr8teMTG9IQj7CZ
ReEbVux1rREUslJPNlLIyqO4Nbq7thViPx72+OdsHjKpFb45dBylevNobnU33/Fc
KC9GloiEwn8gb439QeCWgmI5S4v/hSGRnkLFxMIikTRcPzqc9WCtu5ndhst7jK/s
PvD0pF5Lb/6+6TA/3U+kb5Gto0bpFUUKBalXykUpwav/j90AmYTVqsrCdzWJEN8o
5rWE775kgfetl834M5pGMXpkO8HIXVnzyt6sJJTvPw6Td4zCzW184ZvfK5fgslfl
4E5vxRp/a/hgXEslWFlTlBneEH8mGV1idfXygY/twsujyF64U/F64KCii8dveDc6
P7jD+cIjlx/WUKkqmLzW9UxUmK7q3NHbtJNIHDzRqY6rIwvEYqclwNuxYFPTtNGS
XZxYUyDB0rs1Ja8ZlksiIp3CwsHvFy/o7olI04Xmk8kjTeyAFa964DXzn8mp86m5
GaLDMCDgqc+QIjK7O7uugQlZDDyGE3PQ1V23DHmc6ylG/9ZhGMdgQztfH0FiiPSw
w3mgiT2YQxSlwpC0eE4GG4txqzQmLqedZd7st6MwQ+LVAoOxg5pVAnVSdjNUtFEd
BP9q05PsPwjXSQbVnnN5taDFOmxxmnqzHeMYmeX14WdqJUjj0Uh5y1DBquZSKP1y
tnDixfYAYscJWQ0QNGQw+k6dCIZtcdF9TYEp7XsrzYBsoqL3AehQRzuCP+7KhCQJ
6PHHvGMsSogNdgVJn8V3rQHVxLNg91A8U2DCt1ijlxgug5YzRfoM9/MWe+9b6fM7
rQY28mpL4IhjNJUcvkJj58EqljklLW6vdzjGP6N6ar64z/5QSfCUPJLfe7+HoXxG
vZuQgl8JakEAOFzDsZFdHeTm2B//OAqP2v/5ar0nuISeWI9Fr9jZDqRNSJx8vX9/
jl4FFF8hry/i0fg5sp4nQNYA2ZGmliw19H1otGGC/3wj3V9qZsGgJdE5pkAySA9Z
YsgVX4mSrsC85hIp/oj+DJDJq6BytOOfgVQTgz2NVw6zDToapooR21dE4KyCB7pg
MOfgCeXnVQS0CPXmF3/dFg1zZFpchkPEEYwSwvCZK71qpYiSQO14qKS8lCRdHhOu
KQgBXO5TukajTdoEffSFJz0H7fYW/v7weETNS8kRhupC2f5x79i+/BAQUbCxv9Sg
U6m43CrZCu6Xi0akywPAE2ucVSWPaGFUBOaW9w/I57CUh6V7hB6hEhIia6Ub+6DP
GKs41yvh8VeKBmfkoU/Sh2PQp/bxP6M6w5kJ/jufzlcKWtHWtAckPohqV2MvtYsq
Ewy1QonJYFBHkFSI0rLC2j/vE1nL5ajgbyB2T+KGq+SFjYhP14BLLiYKoqbYZf59
tNUcx/EyEw6l9rpZeL76KqXzJKP+ezeYVtWyNLZB9lAhyPMraeFyiIYMc2Bdrdu/
rYFdBELve/BOUhN8gt222MMLNQl0qUr+W6VDd+xU/5IpUrkNRiia+HDj/OQyBxdO
NrzrlDH6C5ENaZALR4MAfGLndz88szM/doP81KpphZ6FNFBMyT+iNJtE37Qgu1rq
uSXPcJfRd+SJgbP20bmKao5BXvCmX/lSnjKbKpF+ngBLB0ar468Ac6JfLqpzfE3r
5fsK7UhU+61w+x4Wlj8qGWTAway9FWrjmBPJ3npTnkfeD+0mLBTazjl5bc/E0gf7
uxIxyQfby1vgDGIZdTD4pPhbZzpqoH6fkU3PGaUhb0m+Ykzo3d4ewfy4aWRvZiVq
wkppwzEydPTqfE/WHfYIidb9qzeCtrooE5pfxONQLNOtQpPMaqxnjb4IwOfhmCOm
P3EkhFBrBlPWUocEJZxGTWuVdOhHxRzGI+XCNjhrENk/vBeetGsONZ5/uuOBDow6
9UJ07hkEhC+6l1rMVgGzCEuNnsLG56T4/WYOy4bfve7xl4lhXOjlJatkCPhdCfjR
2Qt6GDbbOFq3IVav5VB22+HdmgKfZzl81q06dmz/SwJ5CZXo1V6Ssr45/mN9wQZa
MqdLlZSMw3QqYfmShAILx6wzt3bLXUelM5SsU+dgFEIAcv1bqk+TxSKKi5WA00d4
zssz04DaPs3lV0II8nmBF6agW5+7HRb6XBU/QQo6wWrTNnEuuDbBQh6Xtu4y3PfB
qMXATblWp4+cJXhn7LtJYR0V7FfH7sECDc2lL/jWBij7PE7/S8R9efLCcWzTXvEx
5D9ERqZ14uXLCjDe0pXGz7+OEQLQvNkmE9DW/TXyK2Tc+VMvhPs9nDjTR9EAl1Zk
DLk2CpIt/jGLUKkDNXMKMxM45p0CID4PNqXUDEoWF4ybmfWaQbHqIP6bwUVkICIp
/K6cWroDeXl/HFDbPcLz8Q9xgX0aMG4h92t+zDss7MKXK/Zeymrm6rbaUiPzfSC/
VnxlBkDFEkip9LUHlkMQACJ8eA4zeC9vP0JV8y74SsZm6CZuZV5nx16GL7WXv/Qx
tBUIq39F9BcX7r7/c7TyF8qg8kv0tZLpZ+LzJyoutP7Yvn58ABYY7tP0JBUkaiIH
kMBytsVI7Ph04QT7h7ReXv4tx8fgOEwuFRlgOpdXqPGJhfFp02P60kHdNwopoNcs
mJHnUmL3cgk79J1h0J0CxVG4G63GD6gR+MvjChX7qN3C20Rep1Myth7Il0oSFHOO
iiHe1xjGe+3ZTBdErcYmtSN2a4a5gmaZ7laNDCb3QCR7U9X+wBjegqNdZhhQl3Dj
w6A//Xj2Kzd4p3D/IPAUZ82JSS0wNTt6iAqfbAw2PvFAewUVe3m9Nz7AkjA6hvzG
e6Ft19oSh5dq+zjkYICDFSzMjZbRBQEys4GW+cgf66TeVAWtorDmvLbJB7wKre2v
uf3dZ0dpsxDeq2K/eQKpWYRcCqNegJFR1jOt3UAeexP0AQh6rxUXoFRQ70Hd0FV/
4pq6PfPKKkEmOkvgDSd1thqQrfWWfCXD3BwecohAAJygNphTqoblacqwyLWYSxEz
TnJHv2usZJ06f9O8g3EfGOuMU5CZvrpTO6g6LFj8QWITeLIn4YG+nCpX7mvXRY1w
c2DpVAvr9fszJhIyRM+k53AuYjvdY0YmXLbz31zjqsLBcaGgOGk1z9ZcsqGIjszo
otd+sSTRmUGsRp2mOOo0TFJIvKKKd7c1Qg3T1dRrXJClbOOq3E0KeFlBGsftsRHC
civ7Wh0G4L+SyQz8DPIQVFt/PA1DX2x0ZMZiXMr+/+jHN5HGwhu0AHFVeFZi+BA2
Q4R7g4fhe44TfiPYe01WjHYp7o4lM5Pjmj0h8cVeCzWSRpKc0qmgAVy/hF7vYLHA
D6IHrsK52wt7N2ec78+RWDUaMYFJyWDc8Z/u9Ijkto04LawXMXKvkuUduP/Y7X5E
6Ndzd1KD3BY3rMwL5/4pTH9Uto+nAyv6awGfMeupzLe2m9yIemkNtZv+t2ZyJYap
7913CDFen+1owm+MHVzKxIQbnJgyvrYT+zSnQiZhHqO1xl7vEOVidsW/R8ZA3rHZ
4VA6zIDi8yoMORZVgAIyWonYPgY8UpgpXju1nmTdHatiTxHOxEZeoxu6UZri5wJe
eRh1g+CWGr/l9R1xJ5Wza6LXUZzwwTo0n2Ux34HIJ7tGdPOXZ6W+lJ8IMx9LLJkV
net78+zgFBfkzHjHHZaTxf5rNhrkUCzzPTBRGJz7ZcS6oAkv0YkIaGrQMcw6jobv
+hQIYtbMa2SOZF4w52h+Qeixha3Q+Xrq3oqW/AiSCyIcUH1zhBNJF+4IE7yNxqH0
8dq3EYc4oFJzHYpibNQ+h2davij7lTeVWNYBHN00U9qgjg6KPbpVGefmrcJn66UW
1ixOUVdo8MXwO4UJHJFYv/MQNL8zswO+jTeyhEJFsPNFJTMlmaplmHffw/FOWQge
Z2xuGbaHFPWdg4PCStBvrTCGeKjVDmQ2ge434mvA1lqj+g/AZN4kIoQhCxMQWb2w
QVIqukdmyGbBWfT53BJUKfziQqvjFAexPOgRw41K4hZ76Z5lT4Dj7fuhL09DDpXg
DWNj1n4ij6tSblXYV3EInoTE934gXleeFERooTJ6+loiyaExMKW4lIrCPYE0wfLf
SNB+KltkvOxmJvzby7t3AlcRNiNBXvhEaeI+5nqU0bgQqZZJ9xyFyBUHdxZ9NZ3S
nH3qImbJ2vhWVSEeFsQUo7M9IBcFjOF6ivUfYpV3kjrwRBnOHstIPwwvLCupr3US
F5QeHCeKRl8yEOZYBxP7gq0tcelkZG2LgZ3nRWJH+1wywBuUwHTB2xXb3rIBd3fY
xbB2mv0ZjuuwdUgrPRn2YlUUcOQJ7Vw2JkvndN9XeJILygMozB6hqicQh4YAG935
MX8dQZIZZi3JzOxQRpBn177Seme9kTPP4AznOVmzFNuwciGUAJyQXkjx0ZbDb6/e
GPSdGJXwYVFMV/TeYIjeb5U+1Io4E2onB2RB/176juo+4hpzxrSDfj2TAKDExiy2
p69w2tYgc7HBeW4/HSJ6SjvnaDbSGET8zBraMobjDTLZrNDHa4XBuK8PmyYURaDW
hkSg8FLzA5UcznPG9e30c3ZFh9wLqnLKYpyD1bbk2/I3toZIHxLuChp89XZszFNh
6eR2caqfkZIw8oMsmsfZuL+fjXBEQjcsZhxdVw1ASpUTKkNw4iNp1eMPqrueBlfW
jVFGtg3IlrEybfvu8CDNLWjdqcA9AwioZTOXq+djQUZU0DHvxvIKbCwXsEGVB3O8
Vle8lAuaiI/m5phUEbmGE5IKG5B7HtOfPbQT5Zp9GhpKQYQymOL5+zvoMds8bug2
MVH7azfPvtrh8BeFB+/b7XQZWkwA5rctQzCeFE1aIHQvsYkxlyBWbncl1gkRgvLA
mWawSV0aZ3IkNyF92CmBd8RmYkOZl9goahLeQGtZsYbY6NGjBvnrvdmRdN2kStW4
21ZxAoaM+vNfdACAHLMeUZpd5lSYFOcPHOQ3FNinH90uVPzWhLOpJyRPCBTuR+F9
OObERLmepcBG9IXINb6e3NeWMG7y5QJq86NrsHdpDsMXY/ax4Lywml4aUyVHaNCm
OLNT5RAQ8fsdAplJoCQv54StjpahCwy39L7pMGKQqq1mFlq1XnXmgNtlLKFPwuSp
7PVhMKHL+fm1Vw21T87Bzk0FOl5/nxzKGnASqvTPPPmPX5tG5ioeIh75KeBExeWA
nfwch51IVlmQ/pcWoosohzP32QiAHGoMSLRO0dITAbG7bCrSYe5llqttFg/pVX5u
ZIoKLLYtjrseAqMi4k6K3bN79dQOvvUw4pZNOu/HDThVWinIctEUbmtuHzQXjLCp
eNNb6NuS3/Bm1MjYtWgH3Czyh7k9Haz43N7PQs9WZG/ZDrI8kzD3pjhTkUXeht9T
faMf2qtaFcEFR7SfhsZwNL+BVDzJfnXX1fnVnQdkpr8XI8OPR6BUoMQKDBqdyZv0
IBRExzvOinYxD3jYK1vnDu4+ywgNUPvYHXjyL7oSthRmLa3sm2Gfg9ofTUz1LXXh
e/zKLLRgzYHSchJUpI1nFcpI7bPwPxWtfou5aWin0mhh+PI+ZS4BeUUg3Mow9Mad
N4BJsZp1CeN5qy5uucigtCm3E4Qd6A0gKR2C6LGBIvrS5wxADY2MWPEsyGVlea+S
jx7pD1QpsmTha8ontFgTQPubaCGbhy7+GNlAqAx27/2y/9308/cr+KECKXWCExfy
lY572xlx9uvqaYuZ6K+VNx80Dj5i4ghlSMUMaM2YTvS7oXoQbMkiYYt/XhtQQbqw
mFQf3TferHji1KAuTOlXYG0P1l3mcQ4aOd+uTyamw7RJ8k8IsTbrUrgc/6IasPCR
t4jd1TldpqvGEh8q9qpmBNHJkGYD71QDEZNfsGgS3pOvIzyPDxStJFBxa0dwfz8O
1ET01lT/6c65eBGwxBGTTJvAKw8xLdgi8AEn707iyqFeeRODGDGlkhnrn1BrUdiY
XGCjaUNf1+08jSC81d1qeHIT1JnPqKcfT1LD8Qu/5w/RzGG0rqQAquM0lOgvDKwD
6NDkqL627IYYSS+4FTqWRGUAeWyF3lWT7jftoQY44yJ64vkMnirpNAhdZhrgNFpO
XrXhjtnjn7+ZoPh7Xkp73rsMyCWa+PG3eOr38s/P8XaROZGze2KeKt+snBwPg88e
aJc4s5XybO84VqQ1HGKcEVGU2FDAfIBCTUkLZgbp/GMQLhqdvF1xxDsWoUqoOSjG
iMlGP8fM2UrN/GRya5gzTFq0cIzHmsV9i+Wo6Q/pamXlkTyLcl1pEhr0o1KYJoYA
TTrj2BbRyYBHdhOxVkGKbg2iEkPB6FuZX4w7gdWMUF/IkiUqyhDggWn67AjotQR6
tRH0gFXsZMAEiyOC6x8yLv24bonhSM4AHsklVfzDniWRX9oxCWyAbW5YsdcDcXH6
19pBGQH76zF5rH8i5iYgScc4UO/lEQFSUGdPwHt7YM94Vpj6UxVi6BtTrLj5COQy
YjJBxKewJG8NX2KJrFhcYIT8AzaC5lHMM3b9ZXgdFEjwb660motqcArnuSrFk/cw
+6aly7m0EP6tlVQ6zYUE8QLJKDBQob7JQhraTE8+CopsC8QjMLmK6LkTrpAd2LdI
A/DmOmoz+rdi0JCRU02+JyUQGK/qFFiMEmMQop9nz3otaFUtAc5nH2vQexWRCpCI
UtumiIsKKSTK2Ie0M/CwaDSLZBrSln/MYeDk7YlLIlokZFLoGmzU4o7Cgtx2rx/q
0ncDjsna7bFBrBUUZ7NE1gaQ21YbObWGQzVCQncoEiRf/V5W2Xr6xtFEepzTQFcI
qNCdylMZjzeWPV9OD8BAruxE6+ymdf8OlMRGXlvY+Q6x9iKgONRjcJxeQS7pAy6G
ObiJ7P+gNNy7n0GC69hFA7CgQ6XiHUxqtnnwWVRp1n8dfad8LqfWTuooqFoIWaDh
XVXc1AnvcZKDa/OlMYz/k/r3H2R36kiknWeUDZe8S2Czn+2oKxV5F0JfG3ftVu5R
k5WJzX7ymzFDooHbw6l//71rPASHTejNGtljoBjMzYe9E8oJcNKz/vfA2aMkQVdm
QWAZ6/WOHS2vpM5W+vVjXlcZgvreCOfKkJ2cZQnkAdGlUoUE1y+8uA9hrqchNS3t
Ubuj8DaOv7AnCm705v57reGPC7w8QNQpfd9jG4ikdl8/hff/XAd4COVG472umLfJ
noWUiWHx6Jk0EdyQfceAEvP3qEg0bIHkppNKZzATLvSMeZ2YmstUJrE/x1Ka9m/i
26yXzF93yHWlb664uIp+biA2O9EAEwo6VNJJU24d79uWCm8u9cpPuLPU26pdI08X
ULtErx6CTn1uaHqlgy0vySo1v3fS9f6rEpbPMZVZUP5PUy7BZ2J4pLgsA7X9a6pD
VP7nSykCogdWv5fp62QdP178am7IlzSqa1jmqnmfujgOJBM/KbVRE598QFJtdHp2
yrG3EQQ91ndLJFwU95uuYSnEe6vkGk1QfgMttMVnLanemumkEzT2O3hY+HZsYMek
PCFY3vy79nhxLZtm48R8QzamnnL7t01RkFciwfKnaFmNfM//nWnU5bSWJFCaBq9x
jNTj630bJgEjwJNa1MWSyJBQK9dy70hgteNiIzHcxB054XoZQ0fO0zRsD6GechtA
u3gmyVmTXVL4l1MVoyhCje2XVkh0rXET24Y/R9NaOSbEqyY0yKSo8phpRCLGt+Xq
Yj6XztlmPKOmEMOdG92f4MRLQQ50ey8nDWwp2OJhdGHbIHDlPhPeGJmO/Q7FwbP0
OLz3K5keSXqT7lMMH3JDDXmtU5VpgtzTf5cUvcA/wbJu6Ihq1RAyN1qRvLnYvrD0
jwZD7CCHCqM7a4xLT1kyPGhxr009bdwAH0msXroaJ1GDYYFURzTY4DLgVGVWXG+x
ZK0rJPV0yCUKHikq6UMV4w0Uo4El3haBjVtumpljqoJzc8dlhZn4rP+2BKTEXezQ
dDglIbXrVs4qwV/73004+NfMkp/3akpZbm0fQUq9kbU0TxxJgktKYW2q2PnMITBi
ZYu4UilNlXtk7Ra0jg7VsWtLI2XUzOqecdvOEFyqYyCyGC4hBN3u1wXGkB7uPkc2
1pBiShBFypnzfvNH0hlqFBVl2zBxvXzVc6hUkJqd5Y30mVfn1nn13uJjBFBOrfHn
db7q9tHKBWmtHuoIHdsD8cYimyu8mbHZZY4/joFMcsqSEFRB93EDLG+ICQbqjokM
NO0LpfL3u1gKhJWjG/94KAb6oGZUu0xMgtg6+iKoWuFsT9pEK/hykbR/yPvaNACz
oovRN7gNZeiuKInV6iVavrnqPbVNTKKzLteK2epkkQvmMPMGwNgjKgb16V6gNxa6
NX/uvQfzHp3KhfCjuJByjQzQJ6h/VHiPMc5i0lFHlh4VjNqCgCjeU5Z+0/KI0AOT
+kkqTlVki9uTUsfNMOOFfbBC2mE8UjPtox8SF78hCPkpy4fmMjxhD5dwS8Rv515r
b62M+vahEdCUuHNAUrY/gjo2y0tbFmNBARNCJz8FMklGoDt1IrYToXxKDA1gshwe
drV7F2l3smFIBkjxeYD+n5/uLhcF+efoTBXNQ0XPfYFsdstafWz321aG24KVuyMC
uDQydmALRq2LxhhpwBPGPFNUTKWaVFoU6t4WiaV7aUNcNS21LRMRcHfgamlee/mR
OUNkCA8QkiUghpsrC7o3D+PwStrX5vYVxEBFyWTGDRppRV/JxjhJCha8mMQx/yS4
wMEvRkyIMcm6FiTiPFf61WKTcn/THBU4gkGqubh+cDNX1j8RNi8pgsBDdntebOz3
anVWv9AxXwaWYqZ11Qv6zjID76mjo5Df8MOhvzmZMs/91Jyw5ac0TyZmsYe+5BP8
hnSsJl04D782Q3N694DgnoLeuKsQGZoNdDEFTw4RNbeGarIdACM7eB5xkBGnJIhq
Pqa9oneKoE4WWylp+oJjteP+CR9i6iGcN+a+jFySCjjJ3BvoSrF9tDv4+xeOTgq/
QtCnZblLMDJgZbWIizuZuUgN2YK5HZ513aC0iXO/a1d3XKFpauzXQokDeK1Bt/dd
+ml7Zr1hpkFD0rIGk90xRN2cYkOITzmbiK1ozP5QymTko2r2Z1W5QWkhHSntSgsf
KsIVCalaY8UmMuZKtVuKVamgz2fgSsMg9FW0Y+KQxUU4ugHlVBtEzvPvRktsITIk
x5UeRm1+Haza1fXvulTwbMY+xQvLWHg+EmI71LUmUGVNVXS6ROBW8dNhpNsDu7vh
s6q8fab3629TWc8tkQ63m8a2e1EV5ys1oB3PfwtJxx4tJwqTo9/2QHw2gHzw6CEn
918/32toQ1rGV+4/ZU61plpeI6EWLgANng6cLpa80ba7MrqBHuWkGrN0E0ctyPQq
uhzoSmYrRHQe8eeWzoxfJsnjHJtak5Jr6p9JEjI31SHwxtyUqE8MrR5CkX90GKoE
tCCaigVXaEYL4TomrEuMSWjAUZaB38AcnTuTvsbXQG3PXWSxNyxLjd0Ff7twfWhW
oSBEXEUZZAuAJxucHjR8nrHMhJgmLUUXWfl2jSmAWsifpEuA+FJEI6M9777irDDH
vtRj8kPHLOvBArSESwV1pNY9eAXxUFUUwCOJqrpIqaQkQ/rQ99BuAUZOEIw9bQlp
vYzHkSYqozq107b/yLOp50YxM2i25pfPswr+9Sls0RdNd57pSMFgg1LET0hBmmcg
aB3UtI9Te9y3gTF4VP4v/xbiF0Ul+a7ravhWnVUq9t+oT1kKX/md5NT60gNxj3zG
GovD4Q/QXtTfY+lmFcFuSX95y0r3hNkRTcoZkZOKD1Uwd8jSSr+GkVGdi7xGPN/l
kuytMb+npKxyIOisXLaZ0qQyAj8ssRPXVP7ZRXZLXNxbWVCY3s2Ey4TlmHPr6Iqj
/DpBnfdrwPE1UgOZk5Qiomrw168KCyAX4XpYN5ZD67CcRwNFkICNE3PE6W+Jj69U
mNrcgwsz98feekWm7m+2bi+VS+AXQOD9lJos0isALQtSNje7HQDJj8nZewcWeigd
2L2n1tede5qGor1bkoHvaVXE2//6J40YAkmmvvJNW+DITIl7nZ3OzPzll5K4KAu4
muX9Cr4S578o2PNx7pViFxTBeiDnkoN57ZIDaoC4KXUtTStKkOD0yinv79MHfxn2
aTyAVGXvgPxffm8MlsFC+KEhQx4s7nltz1jO7l2ZtLjYsu1sJgS+vYzBZ0gzRGIs
llhE47KlqI3O3yCjns8OPoHevziJFzo+H9GR1mB9sRp7Xcjp1tcsfNJrvbU6shPA
ELCuUCYRzol/Q+it5nc2kphAH0otRphcg2prgCrgC6b14Q1g24LQjmItPAM2gc/9
uym6rGatj+MLJo+D6LVL1icmag1LBpJz4a1x/WmdZDCP9VIa9v2i1WTLp+cWpfEH
NktqPn3z8WHayqIDtjY3yw==
`pragma protect end_protected

// myPLL.v

// Generated using ACDS version 24.3 212

`timescale 1 ps / 1 ps
module myPLL (
		input  wire  refclk,   //  refclk.clk
		output wire  locked,   //  locked.export
		input  wire  rst,      //   reset.reset
		output wire  outclk_0  // outclk0.clk
	);

	myPLL_altera_iopll_2000_nw63ofi iopll_0 (
		.refclk   (refclk),   //   input,  width = 1,  refclk.clk
		.locked   (locked),   //  output,  width = 1,  locked.export
		.rst      (rst),      //   input,  width = 1,   reset.reset
		.outclk_0 (outclk_0)  //  output,  width = 1, outclk0.clk
	);

endmodule

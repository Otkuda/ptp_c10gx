`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
EnXb6pz3Za1VX5uyUSaesrKKJAB9G/wWezkFsGMVM8YxTqjZLuSmROxiekPFx/G9
SYw58y+OpRZAZWeqEjqtu5KbqnEX3xR518vXbYDF68LBIWHOsrcKhZ4CYpm09vTK
TtA2LrEBAZT1M146KjF6ukUFP5HTJH2CZn6azXJlSXs=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4080), data_block
MDUuGqDkZMMUdH7e+fcjMFYqVclxdnupXWIdABeqz8Dkn9pCqd6RP6aIRx/+G/Ar
hSE9Sj5JLGGzsaoTpPCh/aU6R5ov1JQaIpjx8BlHdwao6E+aqxY7CRwJp1d6WYb3
ssoAc3krAPfY+JcUW6ZfNLIOFcGGXKqL2PqdQxg2WX1yJnvv5I6hIWxsXQ9nvBWs
4nv+U3pTw28E+MlO0c/el4qlWqtp6n5/tCvc5eSyR5xMRT4JKarXRT8TBxGk5WKq
3fmojfDb1Fr1u7Sg+PtCvi9H7RTH6dZzizy1l0F8GmwI45dRC4C/6DYUxQtA8rVU
nVvUQ1B4ZJQm5vuv+WsViDAILH9SIvu/fjSsmyVvXtA1LSXilXQDmnRwuz27EoUl
PODKtoRgf67r7/CRoOLUEPh0701J/Ja/DOW7RWG87CD+jLYVT4DFxYEDCSoq2/XX
p6hv4/vsv97X7EdES2Um3bR1es8tsUsjg8vTUENq0Gmk/3nZbQeIYR8izJAV3164
RENQPQ8uoTGCvtrXbxNB3ewLJk8vS658IiS3lBJj7g/J01/ADe4qlh2SAs2ruE5X
SDwVvB40OtJTyCN5HIpvVgHfN30fpIQYF24z9YP3FOUjvWtfnxM1B9JKL6dmU3yf
51pFyZp4nF3W3rDYTb8K5glUNaQZWytEN2yTsThWp4SkfnouLjaHEERgdy3iPUsQ
XrBebJUrcGj8qr2Wggz6wVBPCCbEWZD0NayXTWGNp2nXXLnlqMO4IdA0rP+ghXXD
gWO88ptmu+Nj74dNwp/lDu0ZMCaCdLGv8noHUTLMIHkNURNdDXax3nwa3W5qRwSy
I1PUtcBNw2E4/MUOOKW3/LLYP7y88bGnNT5d4RnMUy7SnRJa8AyEfYI0aLKbps80
Fi7A0G7POrGUmUWi2FC5tO+6DNZ6GlvbmiaFgEXb7UUsM+yPYk3oSRC8qeJQA8d9
Nb81rfOc2zCzhtgzqPzlpYBgpj3aejKFYzTTPNsxDXBDUSFcs/BCuDbeHFdkonip
3G75KLIRihT0FcQRPYOEyrDiVXiV0U06YULk4FHOanGdc0jBtO8IcgYV8ja3ssHw
mtKBnM8lWnI8I7vSeBlLjvqoMEw6ZDVfYWqENy1VvxZnZRLyp56Pbg//Fe9htKtj
7IIcdu86+TOdn2YEr4SSM5vG+8kjqxMhQoVIXK33rldEXq2XevATEsDE7inofGWJ
6ydzUGksEaGrCOq3ZUljl3xhNBGhRPZ7EEK9zpGIyjLZHMZrUZAxabO5AWpEpo1l
l+oLuFKEFlBjKyOKKUduO1SLsYUgza5B98LoBZDYNsiMPAX2AxOVrmlzLBJ/1P1q
zv+nP8fueI9teKaE6fNP+TYFAIjIbbXwL9lBhBjFPr2mNTFBXjqmyQ9UccNLH1R+
3mmaCF/DvBA5OIQGH9v9xxMx07fSlm2xGAYcm5yUuiicyR05BuSFvpZLNqXtEhFH
zk+QZnWnvlQdKI1PHuv9NaH26m9v0LQNo9/JAZAYrU35utHaXSXIRBuKA7JxyQ2u
OqGH4eAwjeIIooPO92dknrXQqJq269n2x4iPCgkKwYxaX9YcxEjnuGfE19NR9kYT
SBpmxpyhor5vdueiGWh3wXt/lFXciV5bKhTmlT33vrAuEL34dz0Fyu9O3jZsKQ5y
bpdK9/tIMNXGVLseUFzfFoA6u7jS0//EiXOmpRHaVnKZkrKcgWaO9QIR0Ro8cLqC
/vriNlSzReOtF9TcrwpcXOqx0C5XnQ6NkyrYC416s9zjvioXH8vRBbu2bcg6yxOS
ABUs5JRClfeZBS6TQ2rMpStybxfbpYjj8DcnqUO0aC0wknwDyIDE+WqUbyajWvdv
ZLrtRYnfw3ox7h+RQFxQkeGjA1FE4oaXka2NdAIYTLHoNasR/RmjOZO+FqJYWDR4
/u1yw91s+9RkI/EmOlZ2183nunPwpWIzhpFY1oy5DIZBZzgWvYV/a9+5d/csc2br
+sGBEuTeY2+BFIBN/bj+/D6NyeDjq3MtPW6igZYvpvMZJ4GgEvxUXAeNweQ54TES
ecVhNqz1kbJf2Hq0LQtmtij6E5l4xCfu3gj1wN55PZq1Q5roFaQA2sNN4pGJZiYD
XnPkXAEhC2DCOsmE56PPaNHdT4Oxd6MYe2qeScwQR9KVn3Bh6qrThVVaQ/5cIf1m
FvpAdkxJFQuBVmT8XT7QvoS1Bl9NFFhFgWQPVfty6Ggub6joWF87ybPm5uUepTEW
6L/bXkVPO0m6k5HDrG3g24Tz6uXP7UOR70vcOKZ4fDRswqTydCcFTTdFeXA5Tnv5
2axO2IB39iahZZbvMsVPgeHEJ9pextg1GhkoVT1DA8z3nMu80sqyEmrQG6FbII62
mOhga7El1hR1I0IEDDfeDA5O/cLK0WP6NmNmeZWGg0zTYps9cezPs/gNUDOCto3h
X5CPiCsVBfJ037OeSbneNFWwdAZPp5zUaSnz+Mccyc1Yj/sjTMp+K9CjnNQkI45h
C2xDCixfCHj+M3zfabdxfvnvwEwU4mPyRxV9pgIN8wZdJfzwNqQWUhZM/4LlyHnN
Bx0qYam4TfkpbBLdHdXDXP+ousVPIHNQ2xiBDqhgD7v91xxafpVuHiV5eU7GRBLZ
PRgfGdBZZCRUQqI4HPjf/GQsXrc8JuTbmcWTUjgPSrzC798zzuQVNUI7U4ixCmu7
XBHe2z3qGWJWcY/dxyT9pAe44m4GdYOSJcFUuxX9LI33atHHXxXKc4v0sLItds/1
SgHsAbNPi+s4uYeE6AnzFx1hpn6MQMBYNrNeZzQyFPo7jV1SWQdMT3dB9KyNK4G1
oEZYAwN7glnMWEXR0jhVDj2dX0MmHxmVnbwlcsJsO1caIkFTr39jrxtJVAJ6xNKh
cMXPqYX14lGwsL92zyZS6yyMt/wAKaKbIm+lzBZ8klQCccbv4RifuXwmPj3oZ48B
IpgHHn5fV4waBo/VJdGxBMyzWSwdpPR3EW/WO4q3ujta/UfYVFNGcpJxSyU2uVwz
ca2yvTVnN5X1Rm1Hh+U0HsOsom3+1uEcV132i6QI90Dzubmt7ptwdfoeWWo064IX
Vhgxv0HJzPaHdMqNus5/BE+GDn9BHV2e1GPJy83Wx3P2KLAMp/AYY6ql71H5aIf0
KxpOPRnYykke6tc3aaJc1XZk1F095Mjo2RMJ7gXuNqQ7ewjbh2poMmRXegfh/RXE
Bi2rtj8XhlUuuhqQWYn6iJxWG9xzMXaZPLLs/zNm86mpRh9Ng6g96wo07Uok0XRE
zmwWx1j97EzHQjWyEQFnD4ObgOgLuvGsrkWLQ7AO24nz3HGcsc7gHnyuB4UQOw82
21pf6groazCMUHNi0v30tLFLyAQe2TmMF2jnq//i/9va+uKlr9amAvQblh0/17/l
t1GF0ML/SNQ27w9jTQJdjFpBSy+bznEToIfXZqnaIYcGCP6ufsCpeICKJA9ZeBSn
eYS82U15LmmbWlFpmlJ54wzxs755QCjiLZJGuqVT/KUW6I+kwf1THTzbhgbaP9uM
6aY9xCEi8s0ZMF11egH4HqiEHIdlancnBWATysKCccnQIhxujo6MUz1v/MGA4Zlt
3JVn5zcyd3Gyb92MSl0/Gtc6f88NL1+DQcHbnYQOi0Tcf4e2JVdD8mu8ATqy1e4k
we+o9Oq6gyeGGI4MEy4yw7q5yS4tCsFVBwmtpWLw/zKWZMH8HNfJ/+agLrpln0BX
NJ7Y6Kf8WXwF95Ow+mBdLFPx4xS9kQSbaHLvex0UAIkR0GxAIuWeeHoe0HLBccx/
4qWnsWJ5oR5azWeRgGZsUCEn7jb24j9Uw1kDL3hwgBkhWfYxGraUNVNXUbfQkKt7
94giRnpzdlvMyQrKBNBa7eD8Gfo+h3GcHjxfyLaTBCStufP1LYsATNwiOq6MBkqV
avFipSxW21P/oT0ozWdgTzgnhUqyd5cIe+jYjXxEUTz97k4eVLhHVsSz03zcIFoT
cRbxhpeDdkcJXps34G3woM4Cmhvt5eTGNN92hcpOsUJ5742InrzfgFVcPSQtLOpR
QNEKG1WyfSadSp1eQJtT8kP1aGY0pUoklFV2MUPkz0Ypb/tk1acjEtyBZ30zR2ca
6BgcFeXSsZWU2oOH26d8tYUvNXttgb+IkMGbbFfRMTLTisQFEWCG1gV/65eCsU2E
jEALDrPAcpsawm8QBdl3vbTvRye8pDv1w8W5QriC9TUILiOYXCoZbPdcU7BOU8Ki
m15KKbc9+yuytU+Qkva9MlO7spJzkLkkYL5K5Hfr6uiD+azuR/Gx6HJmPbERli0C
/Q/7V83Vr97iVS4gJ6nHB1NEFm74e6LeQ3x6o9lGxN5r3wLIyw3Hp4+s1hp6Cpu0
LRWdnt6mrMpMPoqqxyW9s4OjMwxdpm2kKYh6zQi3TJqXPT5MmWUgLivjgLNJoxyl
KLmblLyim68cuRAnpBOopTMtErvtl7mk/YZvVD1ekg2jszxrzI2/SbkXLzwk6KKd
jZRpzcF71U21QS1yDm3BsP5Avda41ob9gkWN9esiBYwrX8JIquYapF6CfZTSi5gE
NVuudDxryKV5SS+niZzalWYsK+XPOFPi3xsZnjCndkzpjqpUo3OtYL+XrkkH7hpr
/auK0dFiIE7PV4k6a9aj4Zcd3OkyjPHHdgsYZ1+msZmUkgoK5iEBdgrn0YyjKAJ6
xm5DTZGAqgXJzUQW+PfHGxufUeYGfpCOn81e2iz9f6A+hiKe9duSzGfJkWwXz3St
3+Dhvvft6AOXFZev7ROnUcofUAyaXXNcVw+kb6wWyz0piUDhl0H6tItM67QV36jW
CWwrcCZ1iE0f1WB55ZxRRxlF72BDSGoO9SYXo0qKU9Uks5z72A8XBHQT2PsJhK8a
myWokEq6h30Hjvgm4wKskOsUYRYnlDfmqI3UWNTik7WBNeFD2PRtg4mFOVA6uF6c
nVG0u2HZQZMDWzhlZycBAqdF/ik7pSQfnxJtSFI9KdMvGgDcXK4ZQ50QQQ7Wx8eK
/iKxzJ5KWvO8P1VPEvoCWXewpVkE42BAOSHOXw+89VwqM9ZFyvPGWvXMBjfKQGRJ
o6PeBb0UpAacmeM0QDZNdVr+MDWsL1IfwDnZULRJid6P4f8tev12TaY6UJZdBHnh
46gfX0dCzBdJ7Bu/8CfNdq5Ks9d86Wj5uz+8Xkvty1IVowD4WmyX1D++0NTawmRB
NXvg1r4r1S7wyU/po323FOZkA94M4nWWV82OMJdAEP00pyF7CzLYjMbsG9vyqWl6
XZc8d1whwBAJ8J/VLDB4xZVn3Gw0jiAz6crULew6ewh5K6/IS8L4nJlEIgAiounA
ruwke7DMpTjVgPNo3q9vXlc52wF676ygImW83V2FbtUERw1XynMflw5lhiBZOmh/
fsCnbJXgKPbsng+RBJxPsixYbkPDOckpbjqaF6Cqlj7xG0jiTTamiCB6kMLs0XHU
`pragma protect end_protected

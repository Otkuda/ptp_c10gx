// myRAM_ram_1port_intel_mce_2011_f6dnnqq.v

// Generated using ACDS version 24.3 212

`timescale 1 ps / 1 ps
module myRAM_ram_1port_intel_mce_2011_f6dnnqq #(
		parameter SLD_NODE_INFO        = 270036480,
		parameter BYTE_ENABLE_WIDTH    = 4,
		parameter FIFO_SIZE_DELAY      = 5,
		parameter QUEUE_SIZE_WIDTH     = 5,
		parameter LATENCY              = 1,
		parameter WIDTH_WORD           = 32,
		parameter NUMWORDS             = 256,
		parameter WIDTHAD              = 8,
		parameter SHIFT_COUNT_BITS     = 5,
		parameter IS_DATA_IN_RAM       = 1,
		parameter IS_READABLE          = 1,
		parameter BACKPRESSURE_ENABLED = 0,
		parameter FIFO_SIZE            = 16,
		parameter FIFO_SIZE_WIDTH      = 4,
		parameter NODE_NAME_DEC        = 1380011313
	) (
		input  wire        clock0,            //    mm_clk.clk
		output wire        reset_out,         //     reset.reset
		output wire [7:0]  ismce_addr,        // mm_master.address
		output wire [3:0]  ismce_byteena,     //          .byteenable
		output wire [31:0] ismce_wdata,       //          .writedata
		output wire        ismce_wren,        //          .write
		output wire        ismce_rden,        //          .read
		input  wire [31:0] ismce_rdata,       //          .readdata
		input  wire        ismce_waitrequest, //          .waitrequest
		output wire        tck_usr            //   clk_out.clk
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (SLD_NODE_INFO != 270036480)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sld_node_info_check ( .error(1'b1) );
		end
		if (BYTE_ENABLE_WIDTH != 4)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					byte_enable_width_check ( .error(1'b1) );
		end
		if (FIFO_SIZE_DELAY != 5)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					fifo_size_delay_check ( .error(1'b1) );
		end
		if (QUEUE_SIZE_WIDTH != 5)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					queue_size_width_check ( .error(1'b1) );
		end
		if (LATENCY != 1)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					latency_check ( .error(1'b1) );
		end
		if (WIDTH_WORD != 32)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					width_word_check ( .error(1'b1) );
		end
		if (NUMWORDS != 256)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					numwords_check ( .error(1'b1) );
		end
		if (WIDTHAD != 8)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					widthad_check ( .error(1'b1) );
		end
		if (SHIFT_COUNT_BITS != 5)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					shift_count_bits_check ( .error(1'b1) );
		end
		if (IS_DATA_IN_RAM != 1)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					is_data_in_ram_check ( .error(1'b1) );
		end
		if (IS_READABLE != 1)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					is_readable_check ( .error(1'b1) );
		end
		if (BACKPRESSURE_ENABLED != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					backpressure_enabled_check ( .error(1'b1) );
		end
		if (FIFO_SIZE != 16)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					fifo_size_check ( .error(1'b1) );
		end
		if (FIFO_SIZE_WIDTH != 4)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					fifo_size_width_check ( .error(1'b1) );
		end
		if (NODE_NAME_DEC != 1380011313)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					node_name_dec_check ( .error(1'b1) );
		end
	endgenerate

	sim_dummy #(
		.SLD_NODE_INFO        (270036480),
		.BYTE_ENABLE_WIDTH    (4),
		.FIFO_SIZE_DELAY      (5),
		.QUEUE_SIZE_WIDTH     (5),
		.LATENCY              (1),
		.WIDTH_WORD           (32),
		.NUMWORDS             (256),
		.WIDTHAD              (8),
		.SHIFT_COUNT_BITS     (5),
		.IS_DATA_IN_RAM       (1),
		.IS_READABLE          (1),
		.BACKPRESSURE_ENABLED (0),
		.FIFO_SIZE            (16),
		.FIFO_SIZE_WIDTH      (4),
		.NODE_NAME_DEC        (1380011313)
	) intel_mce_inst (
		.clock0            (clock0),            //   input,   width = 1,    mm_clk.clk
		.reset_out         (reset_out),         //  output,   width = 1,     reset.reset
		.ismce_addr        (ismce_addr),        //  output,   width = 8, mm_master.address
		.ismce_byteena     (ismce_byteena),     //  output,   width = 4,          .byteenable
		.ismce_wdata       (ismce_wdata),       //  output,  width = 32,          .writedata
		.ismce_wren        (ismce_wren),        //  output,   width = 1,          .write
		.ismce_rden        (ismce_rden),        //  output,   width = 1,          .read
		.ismce_rdata       (ismce_rdata),       //   input,  width = 32,          .readdata
		.ismce_waitrequest (ismce_waitrequest), //   input,   width = 1,          .waitrequest
		.tck_usr           (tck_usr)            //  output,   width = 1,   clk_out.clk
	);

endmodule

// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


module sim_dummy();
    // This doesn't do anything except keep the tools happy...
endmodule
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9kcW2D0ZgE6z1bX0tET7yCAU4KKrbgGM8d5/OKLwiJPWKWKa9Nlk7jlsXBEQcAP7I1pQ55BpJWv1uzyxAuaYXVevS7CCOGzatkm3HCgBtHg4n8VwWpkE8IgKfLDARN1cWjFF8E887TOjWqaHqF4dHvkbxiCnyEiOzyJbOv956CQQf/zk20bqdkJ/Qh/ZR0n9z4sYTmRtqPD0fbLWXaN4GV8XVRcclNkgo9/iadNLV55xDFL703T1hgVbEqSmZvjdX8lu6ptSpxLZqQFzv2ewjc8PY/Dm2LxFnyFURd54SLfEcEIZse2K7bGlFE+rTf8eJlqnVahwMhbGa28rceO1lw7UcdBNW+MK3vk9X6U13J7Mu7P8EV0TdHHLxa6h6KHXX/+RpSDOfL54eEO2W44bJNDvVPYBlWdBpv1fKYco3M9I7nrn21aucb7ECz4ONkvKgeBhbx/gtZLGL/oYjxaDkdOtx1gdFy8Yr/5SsK4f9EEjLzSOGUxnERvQ3PGe5EH+FhFrnscaQDNI3AieCt7GxlPhQOMoDQRffk2BJNICm2oq+ty1hsIvv1CyIiy/w+JvQYbyiMmb1ved7a/IrEGcPfP3DMWHKMpdG1jnndCpeMyrBDlJHIJNgVjtSMcpH7Z0N06/wdvkMDxJr+H2CuPy/CPJy9fxmBuywljfIKkK58CifwuwwTSGp2gyOo2QpvpFR555cAEWUwruYakPS10priad9DcO6r34cXQh1c32cvvc3sMx1rY80JNR4WSORC6Nam0FSpHdten4AbP2QwkSHyZdLh6mtKttqcwpe7i9UhUF8JXNtowX6FRvA2QBVU1gF7oN/Rua+vParEdNOSpDjxQM0OYAPTfP1FuskBz9CxoL54NXM5DXXSqgQ77OSGkYEvOuL5R1upHAPJ8s5FSA1NSOUvV+zlr/CyhaXoR/dkeIPaIXqlWqfMvZs7mUgDQXSv+mYlazihpj8szd64Jxzvc7yTHfUDQ8G4OdRA3OtdwePOBMtXimy5Ab4ajHOoQ1"
`endif
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
c6HgLNXS368R/T0YN+ZnOzVOmUyzcZ3UqEG9gXikozV1y+81BXh13gtRZ70kSx04
4bAzBX18K7IcUD2QT7j/Is52Fg8cGIXk8/DXvGkRB+LfU5/B2ONByWMQ8gRAmhye
WDeSOaTDj8ZTWxmuJzybkMSlNMI0q/AG2H5TbSrbVPE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5664), data_block
mLLgwwbUSchH+0IaY0FrS2L9hc9CEmt7E5MWIXzN/zE8i9RF2wH6kKEKfVKkcfBu
o22hb0kJxqNS85HFHp48QsN88g6XaKE6NtFPLp0WpyxOd6TZUU0rppZSPe8ViVo0
Z8HGaFgDhU4B8pZaRIcpvSfxHLKRhrko3Za3Q0aXztj4IHlA+kLQWgWa7VXTlWTZ
3QO14sJlPQQNpXphQoWGOD5at0OJNgpS1nudLRopJ+1nTioXr9Y6fc98YGq8CHdx
2Nm6b9IQys8QIqhcYZvUVRyepm33/y11LkwEDK8BlFpgfNoI3nsqubtwpb/q5EG9
J07XgssY1COE9EuMFxOL1TpwfgKy0Y5A3LnY0SbQ2NJxYRLbmvFu4obzBY71UFaN
R7S/eoGn1oQwMVAiA+JDh+33b1BdWMHj7GEnwQ90iGG6yTFUUlUw2WARnZMQBV3O
KlwYnxZFnaJpTK30mXmL9W9Z5yahIIJk0prV7Es6xf018pdo0lDKx6ZfT+kJiVeR
+nIl0Ug31pkxM75JuuZRnV9GODpClkd5hfjNjThaGiFfvBnepT7kfaq7d8OjpcTy
So+Xe+vinaFyNF+tp7sknpZdkYsqY68r+/i9shCNF5yc04wG+wVv+wxJuOJbjU7v
gS2CbtHMEBqPVTdgwxP8lykbcaVy7aWbsbeqZoBSi5ZawnWdXEn2kqmJVP7tGCMo
Blt14Q8CDFAJk/BumlUPAyKQoo6fBTBmBkkGYV00dvuoEPdsRjNJsxsF+AWH7Uji
vF1+7IdWo2fIkp/zU1IbzC8K7FcOHA1DNP6LI2Cr3znlB2eBa8wS+YXtcq8nBgrU
f4BFSkGNtPF7YeFF+Loouh7aXRfSk7AMxQEDN611yf9lbDgSaBaYUFBrcm+c7Tg2
CRKA+/qwCx4IGTzI4loZCsakP7L24Ti64cskzmv3fL9VVgu4MEeAxS2O9Fcqmjad
qKbuVIgOqbJfVQWutnLnVCrtyL7eykkW8afOVrwWE6i2cX7/Dk8mZPv174PCkyOw
trxL8DBqW6tPPqwId5nPC7+aITjy2DtCmwMslXGqNRrzaqPwttdTRKVAXL4TmPut
NHDIu9Kgafn1pAChHyRaMidmPD+iYcjs4Zv6GOGgQYFuWJSUDYb/MAF6Pa+EOlIm
dC8r/91J2kW3AwHwymjSMKYcWd/jd8MEQLqw7dmhgO5X/H5Te2ohimScUgFM2fM1
SMjruzSzS/AuNps+WTkH/KdQ1K47szCI9yOdMLekWIRz5S+lLrYuxvZ39C25Y1NJ
kn0vXmW+3MJk1HH9AtxzWk8KrzKRobWR9vGee++xfNKpBRzi8uGf+//pSzhdAVHw
j6lP3to1ZL/hatkw37C8Zw0+33vYUrRQbNZPWnNkqbhmUalQf1Tl1liCrtR4Y3UA
nuKlWkR5IviXV4Ahy5hlAoh+3241SHNmDXC9+Om8Ha30BeHUlXC5hw/HKvWeyZow
86CeDfi6YFPSLpPRzH2we9nHMCqfI7cMPRhrEaS1gq7eKzSFlgOHgApav5s47u6o
MOXG4nqEz5f/12S7q/sN5YIjMdmaN/GvGVoi/U1PEGeJhgSvhmTjBnPsdrbQ3jYg
dBNDQUJOg7rsxZyZO3y5jIOChcgbbB4UNq5Exec8oaaxZ+4rsUXvHW/iiEyUXN/B
6S7ov6+OjcodyyltD9XlCiSoHPq4vvHjMVXtwEPefKw3cwYwlgyoUAYp0F70fLdZ
0Wh/iPfySibnjsoEQx/rARsdJic2kJsP5uB/Fq4XLdQniLfUcoSswU005hrHZeyS
9eBiQKEK9SHzr8kBpOU164spd5zHNi1OWnGbfVtdjWDIiBaXj3ljSR8JYG5mVhr4
zg2VdDcC6KCuQlDEN6rjOjtv9zGX43Yk++px9oLSSa+mcSqZiJ/Txk7a455SOVpN
9eZQ5kBUQzmQbsTfmQmRr93GtX8S0ixaiYME6JmudIhhUnQqWNEE/D3bfQM9346t
GTXuJleewYqSrvZnFCz6WyQq+SS0BeARCzmZrShL/A3ncNkVxDkdGhLm9mS42BRV
EAbunePMbsD6nl1UvENL52/flkZ26FaexQ6DfeFNVw+2Lnq/2bJKXqR8qHtPizC1
nrLDGM+xCFV7ZMEbAJrvoV6g0uWPPxk53tVp9a37nGkGICmd95wgIJs9bZqJ5SKR
GsipQYzLuk1zjcZZCmf4sjQMz4uw16bI+J/0MzkpY4HmHxA/Vof66gFVDOUV30A0
hHh21pQ0Vr0AvKEAs1RVYxO7/+rmOJLoyKQPbZD/UpmV4B17GApW0ANntUgN78uB
MP1I+M8mVB5csKVGFaSrMzEu8m6TNhqsrLldDUgSQNRK03lrUga1S60AjeWDiwa9
OZJW6HYa7mCTj3Wktbpu0rgsOQrLEBu0uOuT2hRFmwdbbhzaAWpP1bDhEvuGAtE8
lfdu9hYNjN+0bhkxJFrFEa/WLT5cgofZOXWSuoUvg9LkCKXu8jGebzts5p/RLmBr
U1Q/tBQ35EWDRp8J6qXqcdMgIuVh2jPq/H5swNKlxUmVZdAzu++DRdA342DQXXve
ua/9L6n11KMnveUmCZ53NHCxTFffmfo9qBLW3dkfJcBPwnd+XyYWA5j4YcMOEGIk
ONnqZvT26PmRRNlKbNgYpk00J6gw92UaaPUMdxOGfd7AQYiZfxPjHLWmZvfGm2AP
22pMhmGxkG6UZzIsDwZJBrgtJoJI/aMltSi7oSmWvgvDh2oRz4e46Mj5lVuevoet
/rrtZUtL0ORUHxXB4BFe/5AXa5irlBC42LgXmfoSkVoAm+uJDMkps2/J491CEXpf
1TE8Cn5EmSCxgTBGWQwuGSmHT9iQLYdRo2FKQ9hawziWlq326V8dKxfV+lppen0n
lqLYLfTW4kWCKRIqJK+v7Kazi7Xv5nUbuJimfuLpG58LxfpSm/xIQCxskBUXAw1U
kn/pa+Ovba8DLWfvOpkgzC+yr5m0f4KfEDNYgX15XEWZ5tOBHMegNx5W53v+k1mC
K1iAlQsslvDn7rpHiDKavP4NeAeilubtI14NKUH/ZrtMp8MUzk/Ezhj2JSdu938a
qCCN5tRm53hRENPa/Uetfk0WUlqye9fEeelKSgl7dediv+mOnn50qpQqUryT6u86
fU+CJCJkg2JB9VseOWm5/wEQ42vf0dGAV5skTzjoKcqOMI3xLamTdlR/sBn9USTI
l6tQNM7dXdP7/rbkS9qhhDFrzeHCimd3jSrb3MvBx7suibxWK3ja5/sMHDAlEBvZ
2HqFnvuURxXnm82OjP3+ryuDSNYiE6HUj7NWb1CId+Ziisma20H/T7Na97w93FK9
mFaHrgxVDffBCZjHFz6NuDpihY5mSwUXWcZ4lJENDgx5mCyw2Do2ZKoBz7wBAxxL
0isu+aG4KFRAXvE5SEcTNM+vqW/MFkqsccEh5dc50ZcXjLA/X3nrGaiBfk1KTkTR
DCcmhQdnG55v+s5F1dzHH/GC6IQv+Of7dIl5usgWIvmmDg9ydQIOeRWdYQTf+fPv
nhiqjyaFB56/d2yySB6EmqthfJ84PWpfL4E4DVFT/ylr4gnEc2z0W+5D55DNUnyM
YjYMq7Q/bFiz8JRMBgUHflzyNIPHOQ98rp3tx9fo+04O8g5Jw8BoLeYexl5a1FDr
KCqT5GjXn6DC0xYo5GZ+3v3IJOemcoSIctumhqtfUBDTTR7A1DGsrZQUONs5YphN
P07a2OWh5N2QMCJl/KEP4as90nurCpbykMmh5vLeAlQDy7MNaKSf7gPZVN1cT6Q/
yT59vvqObiva3RjojmZ7NcQ7FyPZlCFQ77qQ3pM2U3/kUnD5e5y7Wzci2lJu1+98
2QjduVQLf9uYapeUxY/jIobEM9Zgoxe+sAOU2AavFFPDhUBI7qYGbXzeXixyX7Ik
69329Lh0NMA0G7UBkWK1QRrHUCURHHXg0RRMuXA05OqrmSw8R0+l27p/5CsSXQzc
tGCoNxix2XRlD2N4bprSSnkUUxIRcDpGkuqVhEEEcmwMSijJKrIGePLxSPOXP8NJ
jYgl1yM65BAhtV7obFpmtr5NnljGPbT4Eg0RpUT9NQpV4EJN47ClHShkMHfg/l5V
AB4mSqhBTJYIz+sOarSHmxXOYFu8Z4yXc49yChYP+dA6G2awfLVJzjup3Tqw7rC+
9i9JICUDlexFn3PI5NxFoxUWya385lCgJHpNmNYWsBWVmuPqW8rCuDA9v1iwKZXO
JaKmog62v0/1uwsFMDwu+WcEYodUU0gPPBbsXm9w/Kym8crq6g1h3nlhuD7tvdOO
iA79U/PlVk2fHG6M2bvqh3GqJVoUzfVKpx33Xoq8qv+nI3KakAP5sRlcMRNkXad+
O29V3jTwEr2AalEg+5Siqe8KCm1VGI+htdFL+hykg/2G9UhkEKbi9B37mlIaR8hL
scI74JLpvA/NLeEsRgYmLAq5SBE7aBDeSZOcfqf3vahQqs4a4yBt2V+gBA2Tjb7N
nNZfEJ0rZCEwFL2FAc1SSWi970cdVAFi3DcNW26MsjzULIwfdx7PBYsGqe2PJyGL
0sI51EuofHZj5nOlUiszy5CG5Z9pk2JhSf0RRF2Xs+0GrItvEvhlr3cNGhB92JYv
dHdeVM1kPMeYsGXIbslTBswL9pLMny5AZwcDSj8+hOQ7Roqu71mTDmwYhmcDqm02
ia5HmVCXTD2KywZy4wQbn/P8harNZRBry0Sgl9rlz+9PEwJ21HiqIOeWYvvV1yvp
AbcEFSjmAliMZCuIqGfwsuOUvQDj8Tq6ctjunN7SuAola0TvKneIAJ9Bc1AVduLk
PlHTpL6u5dwZucuYt7gdKkcFuA+DDUpoDd1F1aLookwPeDDexczPky/2KSp/fsfH
nbMAukPAYo4vD0vwDNZqAf3r0DK9qv+c79pEPB7d9+EhH8/nuxyngAIue/b1u2lv
5Nnp+962/1cR0rC7fvf69UK3yIsimmw68Uw71G+4gpXoy5xTAanw9OOnXPYWa1yx
OW8ROslo/OoJqcfnJ4Ytr1Lsl++vBM+HlUkddHiDlH/+QFWi5/I4SWuzu0vHjk0X
syvJVMY55jT1GParq9jWn95fc7z6FPCfRa5T4KOQc6DSiNgoneHJPwKFvZKw+Lbz
sINXRjHw2Yb/Gt224YEMxXaM9eVODQ/JPwXWlDxq71kwjp7itR9kadV3Zemb4t2M
08D0n5oqH/ow5QFf5ymVKnpjfPeXOZweOXKyMSdHr0KzYJPtJM10UgRiZ358MihY
ecUiF76zuAcTYstd84vzl+yz2N+/uRWG9qha3U5GZJG6z2lCTUHhurvblpfPRVU2
3dnz8In9t0kHWWHdfupv/0nkOeDUgPuWea5UTSyek3n0O916aLJDehynLdV59pMp
C9MlZI7u/tag7uS1YcMffrHwIiQ0wnohJsfV8nHUHEpBFoezHR2vCNB1w8CVxhsU
ZBXpu9YRoySlRQJFEbf//7tiBdvIXymDfqjHiin8YvTRMh/Q59gHVkCpffHskzEQ
CRrrJuaHpfB9dW1aSXPPiV9UfmFpVkgfMu7ziDcJxfv5nNPX6eR/dNwVO/Wtdraq
coTDKpQUDE/VdLlwIiynujz4Poq9giI1uToroO51YRcZhO1ReT8gkl6qruKBMYsx
U6FywXfeP3sC6TF6o/znKukd8ZAi5KzyXidUlBMKnPDC1zc/La58qxHap2Ajlncn
tEK0jGRMS2gTUISpuv0w/TDVNChJqCoGlqRDWzpHcRLWVhdWaBKwlnEgotZPhukm
XEIoWupO1PNY+vj2NsGQ4UFCKL/8iGCVMxMBTsH0+J1a5rmZAUgu2+KzcRc4ey+3
zmYAdqnoJd9tPk3jlsZH4CV/vOkeDsPmDni2QssZDSFj3Z1+rpC1/B5udOabPI7+
fBlMpylIi6zZ8h5SFUHWvQtFNbOH4K60BEb0Hs8Y/bu8driiqy3PLvQ1Tnql+fdK
qVZZuiAiZj1PHgFKU0x7wTS5qtERjFnjXQBlw8jUnfpqED9IIzPaU9Ux7WmAgEUx
9ktRrCaWyY6P2OtPz/uC9wer+RsATx0MfZ5L6xc4XK5BYNj3L2+y8V713hBjJ3bo
Jj/HJlAcNAgvJ56Xji/s9f+8L/bbbUf4owGYh4Frfely/ZDC5JwwiCznUWJMhZ3d
97LexLBwzzQeENhB75Mz3nK8sZDASIWIB+QwVxvG4MrKwgDroRe9q9N2SiPCeIXI
+j2WYPXLbkaXR/B6JSCVFCgyKsZFn4UgNLkUxUeA8CBKJszB3zMV8JdoSazg8T1P
o0vh89r1G7C6TXk6jHG3YlWHfvlkTvtCDrKLie3l4nkb2nRW64StsG4KgxwV5mKB
KilvgpaVi6Q+LsL4X8wK891CTI1rWbbetOJJ0OC7eAbVQIcJPzQBZm40jf+vVJv8
UFg291jkgyAsOZ1AWzJ4yP5R6M//CqaIW84DAJWm/YlJ47LhiwDrFZwadMAAxYgD
BlrbnSIn0iiwwzDburDFJSXAiDBVVkGEHXMoj2eWi8hxBpzukbQ9sjAWUyGPiR2m
0sviLnfcf1NphIAzqQ6I08UncNXxGBFipo+KNcoFU8qnIz9CTLRQQ6TH+sehjgrw
npVv6e6XOF4eYVGmammylUqoUGbrHqNXklBNeEOuORjPpOHLYQyDkMf0XXexjySO
DbAnW7neQ+36xZEHpTlEr/I7tSYqZW0KMaYJPdtpjGqGq0vkpKvL/5YXJMaGxRN3
Y+jJ6rbfhRa9VwxJ4wMqADov+mqir1r7wQPWClQxDBhHG743SxJq7L3Khd/u0whT
T9CZyM6yD2yfvxp+JN1ads6ZSezvh3oLhiO400+JhoQzmvkywAMBTOJQx308q73x
TmUa+bKBMqU0ZXI+uGcTXUT2JDgMz1Fc+z0g+rsWwZhwAEQxXQxQFIpjSIQRp9Rx
EhGWTnIUN+wOmDUYVZOqqBZ9PHp7ngU1DFkV1OKEzDumUvkUQDM1AIQGd9K4oWai
bHi3ZxMQ0+dy/Rl7rBrzjbbaCvlueYmb9oJgPhJOIzOpC5SM0xkgHIjMHSyP9hY2
FOelWJdxiZxiL2JZniFrpZr+A9T/6lCm/Zmj6dDrKfNS6pwpR1mCHLOcjhYWKj++
Kcuo+4N3fDkzdOAqtwGvCHMpCZmtA+O7qGddKwhUA7ePXB0qEHlFfj/mR2gZcpO7
B9WDELb9aYWO7qlDbjui4Xm9iZ4wXKEL+sxHr7WePhc3KR9HeE+uXbYx3seQD4N6
VXvdwyMFCbAsMvITLyxjhfSwoi8S8+u7zC3VNKvzw/JFzUgliNiXIFe7WUTIZHxD
1u6gehKBnmH6kTlvr0Oehh4W3w5j/elsq4colF3FWyAkJuLsd/99ByGNuEZ5UD10
tSd7j+qSQ8EsF12iaGtCtpulyxorZ4nMH/dggyNGRY8qqfa5V2QLsd7/Ay8cN0ju
ELMrOTRCgZ5WopADwcqUDNgIF1vafhd2Ygf3KZntGMYZHHWDw7N8iBBHArraBRLf
+WzL0HOOqAgfWHPjiyuAcDbgsAgIXwip9DnOlzvzm1fEr8MemGoV6YuiPItzRcCo
`pragma protect end_protected

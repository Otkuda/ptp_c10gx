`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
rz9LEJihVqi+b/VgKXGGrIaMWpnVqCCTTdIHpPDAGcve0PB2T1Aiql5kN5mZiskD
DmOUfXu/UKMXxVohetHR39vrBY6F0UKv9/nm4P8BQF+xmbL+W2k27ESffwwlWWqh
v7mwfQxITYShHG5l0MciII0ZH/+mHEE9I02Gvy+wKks=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 34464), data_block
HqSFgsHM2Jo2WpsdbcuniVbaCeawV5Agww7fhZizDe70qP+wbPq+BfCah0wwnEhg
Xo3ldxB0PIjCkFOYPrXtNpQOVA9apOfCUdCLUqBhhJzVl/NhsS/kobUB2ZeGIeH8
wFaEncadstWG4tXT4j2nU7zSdT6s+Fo9sC77tBNgvEK1EjX/04yHk7wKBDLGBHqf
ROs9D9GFVu/DX4eDUcn4s6Z1BMI01XE1wTGyhc7nbygjYz2vDhyQzXyDot5MX8KJ
EYhnn0HtuJlvB//NzEBLpD99IBxEK+yZDeSwIAtKEYRYuz7cN1Pj2spio2309IOo
RdPtwG8Gb5JHCPCN9JWutdLlcStqZ4CINbS2Swng030guxfIJlJegCL+cI6G+BPW
dvkpDDMsTfCMx01EUMSpHtHsYIQqKB+sZndKUvxa9o8GBm3OHZVeilNwvdRaa0az
z4xtaUHoyqMPx7SbDKupT5Xq9bWTaCjYuYzT/mXMgLp5otrLPYpZaC0d8gf2TJto
eev1xuEZ9whvyZMgv8odlxplKC+nIObZOp0WHvoTnMVjWJ/LyjpC0VBT+OUnCYyS
se5iWGbN6UZzsVlFnVGGf1mV+YMKhJQRXormORAy+WkHupKhuULiJAsG8TLvWyO2
xEkumQS4jCWKIhc22+mvfMxpIXvZ0GzcxIL8s+jImJSiLuyySiHMuPmFMRCFlenZ
4HvkoP+y1hPIZkINzYM/pXd01ctVTWapaMtYFa/OTy+1+xJ/quVGwdJG5G+SuvGL
OvvGkj6n5UXiuw6ZY8ILx7pHVXOGeEQG5wN7vJnovwe26McHhRg+2AoZLl6eLAO2
ytXCufYA/7Ihb9LWktjNdNBVIQuAGZbLh1pEnD8mtCGjviIyw2mK0NySb2c7qxju
q6xrPx59uvHznNLS8wfWL3pG7kV4JYEmnNDR7DJse5ECUjf+YQ+rHUHV5xApNNem
BKgv9WzXH0LqkObbIQYu8Xxv5gNWV73HzYAC5tDT+bIvxaYK1I06hv76ZdqdFSPS
v3hqCjUnQm0MeNR7iYNAnM1xzX8MX1djEC+0ouzAkOpE/DpIxqg/CAM1phC1AVCI
xcPht5P0afdyopBUzgifaTqnl4oowlw7QCpbH/Z8HLzW8SptCgIMrIo8Ig13eCSD
vPeYHQjD4D6RPPRr0Fj5x/sIQ2h7y3VrL/OEYAQoVszhuw7CHurn0MGVj3uPfUny
guxUXqoiW9V9kZmeCWnQB++VCRIBMRxoeXnxPTti0DGqPVr3mVoudo8CjC0d1KkA
1jTT2V94tIEyVi85cYxL/wspaK9Y+152qKMiGMIpBPa0H/F6u/wEwo2BRNUKIPzz
p1jZIBN6Afv6ojjPWT1mAkebm0xMbAov5wOfOxNmovOwAL+uVa8SW364ngLA5I/e
g9Y3k/bvyntQqjW32ul59CUowuC59EeWDkIA+B2sxXIyghty0w6t6cr2BSfbN0vx
dzCM14Ux2Pqj9VGW4fyO684uQfCr+6XMUrq+GNExiiStoV8PsGgOjBbITLHEKt2C
V/cXfonwZ0yB6+ZFVtloYOCIQYLYtYJ30+N2XKhPbAsKROaL/M9PEmXuBuIGHeWG
KFYMdcxBLvpaKsS2yKmIb+Gg9oownpQIVAuBESeHBlm8Pt/1b88tidpks4244Sup
jexyIG61Hkel36CDtpwkE3vlrR82BxE+V5EAK2L0lfkT3XQNFAbEQCO9alE0UOXC
hqtiaFB8gVAizoXv/4nRGN+15VJpwHIAlmMpsQiBzH7KYQP0pUmZKk7jGdcI+ynp
bzqEIIAnJ8AxIhylAEMCD4xGLsZ2im8m6RWbsBJNj3YhheDQIvUD2nthLvOvQYpZ
miVMssp0dHkJ/Jbr4F5+P5dd9zdzzeL0g3nbSWCpEFLCxNXQeycT9Dk+Vc0Sfn7Q
AEY6ofxoyU+/d67/cGcGkZTDb6Pvqmb3DVlFM/U3oLTpnhFrg93Ma/aKPWhFLrAV
QzCj4gtufF3d1SXEWFbG9h5pIztPtWAqunBRi27YhjG+1unciXEDtD/efwKt4RdU
ySvusJFlQAnRRhJ+2VfLSFskrh5CQrQAUicSmUEZEQklTWkfK47Nf7y939VNNxrp
zZwjxsFhYkkFagVHmzM05tno4X22GxWsfsD9mcAtWkrza3eQFCPtKy1hdjPrnD7b
rL/2OQSBhNYbl1fZUE/RW9kQ9H+R2W4XfjBGmZhIyX0uP22RJvaFfkMNN2f+cXQU
TCk3DkU66jQ77UpN5opknAX1s3nonL98cf9oa9tyqp393MVeC/hCqAzUhl3u7aR9
Q76ScuC7r61AtxO678lqXOyoNPfgZFHHAErBxO0dD15luwTEEV7NRraWGx/bzD5j
jHhNbabiNqR3EPbL0YuBiE6f74H7lnjAvPwTc61rn6SBsunDaQ/oz/5AFr4ppFrZ
sbYPPmJR7055/xpAfQWW2Jr2WkpsLZFoS1fmrLsUuTM4+c6r/m2EIvheQnuNdG/8
rTtvMq39fZH3rUL5Pkt5LuQq+8mEH1jfdDybAEpO2DP5XdQx4MR4HqBd7yFNXZI9
KH4pP1q/OnQHedIzYAG3sgsxthBrKzDBrOKpA+mtuDHHdRtZ7XhOKZRA6kHHKR3X
m6gMkJwLaHA8N2qmpEmRskevfRAoXvit8og5BmKPPLK8zdrS5zToUnr6Q7UYrDm9
L+ksF1I+csVyGPBjXyd8VG6unTCWbAQwjkINnhyjVqIIZdrpZcg4eiTaLzvDYl94
xqk0h1RkjhswSFvKTgDflUGqBVf8ZnCqo7NWhGV7HxOZyHzBu9ZnWebeFGsGdIgW
rMRB+sPcCvDMGSCZuLMWW6SSQj9oqyjjPjKLQZAO4r1cTol0v8l6om+39cUhO31g
ug2xM51kN1t3S7KFI3LUeizNAgqBgXEKyxfjriEyHO4BmLssMl0p+A53c4AwIn1L
FIgjNWAOivl85iN3H82PTDlf7ln9RdStlEM1O2w3yer5zLKW7sArwnmbNT2mUzXD
MOtIvEios1WVjD2hPwkcqDUCZYXs24D9vyn1HBs+ANVAqU1+MjgYYaPY/Hl5MwtW
M1Ofs0Q7CLoKp63W4fxmtcpyvvYLreDSIU26Ya/0hLIMzYrIZIXHGRl4eAIOtRLv
frOsFtQH2uYIDjmVvvWtsFsNw8ydOKxTOWDMNH/eblHAxBOSR1Ba0OWZ0yzGjr8C
b0hZIu9DDuiyQLUpBlvaEoIbVeEuhOqZW9+ZpvHACIyw4V+ifbVao17mHSWzxX51
RymOh19onCxtMNwfmaGkSyjPs5njxjQGU88JsebX1JNlCSPEjupdNj9Hjvt/qb8y
YMSvt/1uJBEs8p5/c+aIg493algznb3a5xrwCAz/5srXtPcmyG9HHHjFBGvFAnBt
KBP0Tg8Y9uorTv1XjfM8CKgVRQpnmaEhksJO6ODE1gBgS5W85I6jWyxCauR75arB
10US+rNz0SSpqTZN1X9xUqpsdr8riCDihKa2YeOxZ1v09bKQ1BxFYxm2wRde20rw
1RPVMjR5OQOliA9o0H+7mhmfp83F/Tjtr2RcjJNB4NxadedNi54ezvQDRz4CJ0Ai
B0sil0LR2uj5gAui4J0TaJxpj4wqI1Adg3cAFxUMi91LEBcSd1+IKdNnvmOOuGk3
ioE9msRpZwQHBAQwcWUNRQqs77ONmgF6oxO6PkstydK2Pn0fQZcaemnJXyZKQH/A
L7w/16TN6pcsvUbURk8IdWuxLVAlUfnH6kLeBTwLCScRDA4ybLL+NMHet75uzvn2
KDuuHuwVWG62RnBelKYujkHOEm+QsMI02fanYqx65s5uqtFmLbV7x7CEpXyfbHy8
WjryJzBHZqolV3HF1F9hGgLpE+3yWqPPLNCpgiIxBeWe9xJoF2yzkLWf1k8aHNUF
SDj7kk7XZcwgXGIsnd/liG28x+wULe5Yg5EYh2c7Gh+FVd4SRyo5J14Ofvo3eb9A
UjzQU69e6gkEy0i7d8ej+SjsW6cYPSDXmmLOioNkiZq7d6ytAmsDW1hx9pTt9txN
pH2x6X8+1o3yN9nVIf7i/kCeWRYlBzQ53+uxGrxC6WaJwp1caR2DGqnV2fnsLU45
J2NH64kE8L3SqzMRN0kgEfs7GhmxujkjVX/lkjwGw6FcV/cTLrTSBcs+gwCQsX7D
Mh/TZM+OdNh66j2+b1W9GF9iNhGqcBp5an/KPt/0NuVLEzb06wpEGIWAs43w9NGd
Van+PpMcAXrNbk6+VX+fFt0KeD4UqU868/WA2wtanKULuVM9FefK8UgsHrCeRCN3
DumCnyihrXjTOGXeYkDjVLijz0D/w+jTtEOGaOGxq5v/TNM03o6d5DLx0NLCyRUz
AHtNdDB7mll7ep+NaGsIo5JzCEZ/NVq2Jb0SshpujTOiGIVn+38ZTQCJk5w2861j
RurdrJRBTWmNwNRkC6aTdMNS/hOZtYWrJGGjO2YIPOwfPFDRQ4g7CdSBWwrIxwTG
T+QjU1AxiTYaHcfe70lJlSd6ZMYcIXDAlynRXw/z7ZOMnpQTJ+q4KzSrNRoWjgcC
Fz5ud99l9RsJhGDVQPijbJz5WEDz/nPZapKTC7d7S5nPuyz2uaiPfzHjeKRYiuPE
j/i6P6Yj4/VFh2Dtz+jz7hqRraNDm9dBH3JvhDNAtrD/ah7xi0BQvx+r94cs5SrN
xG0IapcfxDDq65KkXDetvEPRmwTJXZV7tzZW9wNKYVPyTCRVMp7KbNCTDJUMeI4W
ocKR+SeUVmZh3A3DEntJX9c/udTRt8ufUDzedugiG2qHAX04qikc0grbaVAr/eDI
0EuA5qEXIUctdEa+k8W1DEe9MBVMBmoipEtakMhZrluJt5j4kleh/xMWBfoIanOo
GrB5L0rksaUewNcRnVcIY5nvEzDXZiCe0yI8xvwJiDyhZZ4NMDq+mXR+YiQhWI8o
A4VtOCNh9Y6222Kp9BTTie6hQrDpruB7aaohOusA7rLTjXynJFKWGa7Nzfj/Me3s
mqlVQmvI2YqRzAiT/RwKBONCAvU7/UKpd0yI944AdZ1YCWVAyAcg8bbZ2JeaESGN
gK3oq+dzT0KMKSK5FCuyGWhbFvAra/JYdcF8Ch7jGPSgk1vUc2kL8OL8sJeLhZZe
H+57Cf+DbQCRwneKw6ePOJqNZ6AkxlxGMDVwi2U/tjAyKaibCHZ8oUB0ghB3NzvI
UEk2U70SB7HcQaXi2HoSsQsA70kyuh/dEMmGqOxL7Y3kDWUW/KvrwwZ93Hfr1Cn6
Mdp1CpGpkNYGrxc5PDjS3o7AOIteO8KmBuWjWEcFvX2mgociZwTajoKZTXz4NZ97
R1IifXlDJA+TPHVmYV51n8VHH+4AAoBKbD2GzRXWCXilCmvY6W/GZu7NMII122gh
ucixsvhRfIoqcF3ivDtVNj6SG4cTUg1xRVCQ/7tOO9LLZfI3lPW+/cp2wL4UtDlB
sGETAKnvEpMO2Q8TXvN4a3Xl4qppT3Y4TQ4yRVQXnIxCJmAM2yS9yePw8+ie+Vug
daMrbhDGlcARyxjd4COf97+eRMAtpmV+BU0M4U95OlP5blpwZUxgXGivP5vav3DH
J9NA45jd5+WSrHGt3DjfrlQFDTVa0YdytnGNbOF8+gzQpPlOC894qO0prOz2ZGQw
5+/ctwwRth3kSzAcEAFHA3tdf/0e7Xo31jMJUaoSC/YLejPMt9BVGZGsuLqaAzN2
QZagAexM5ZBIqYct118/AnBscq3A2mpy7lHYR0W0BWZQSzV4UM5zcMtvjxNcvXAt
rl/gZjCla6B8NrOG3lXSLeXzqsWk+toflnpuW1UT66/Kpx7xnoE8S9C1Tyk38J9n
pEmRZlvZmfZjqR+FUIEF6P3R6S/lOI+Kf6j0mFpRlWtlZWgFYENrOB+PaF6NoZCD
uyeLTNXSUBR371n2fjm2/Ia/FPGpAaAZu17zVSqNEwBFU3u06ygy9VJbK2Cq1vq1
9uWXCNF4EyyBUHLOOpwUKDTfyhyUnQPSQ86cOO6pJ7df5SwT1ahZs9KhtYp/8vn+
cQC28a6cwD1XoztoNx9wCAjxfGPrw+1+YvV66cgCBoq7B9ltnooBI5zPqx7jbhfz
IkTQV/ybr+C7AdRdUEdIawdSpufHG8SyQUmK5p0COdfdZOEKVD0gY10CvwB4Lqfk
pO0T1yB8IoYng+6mGZFsQqypA9zEsdncpbvLzRlUy10S+fcMmIKO72jii+MS4/dF
3CTLsF2N3mkugUJA24GIQWzYK7K9D4zRL6ZYeZyj5ThzJLmlTAuidNlpHD0zgNEN
jz4ZM5Vd3Ez4x2Xdmqn4Uszx8B/ZwChRFnA7pFw1zYhX30QNcC+uSlCEYWi+U796
5gMv5F4O4YDbiFk8qmqudz8cGxRVO73hNM021uucfV43CjH1gmm0Q9i0apqSP7cr
OfTj9F712psn1kVRGaoJD8DwRSHpF7U7lrrsgskmI+wNhWsfEYbJHcGxeug6g27q
eivl2HNi7+X5Z6X5ZCCHXa/jEFHj45cFjs33GpGla3dIgLqGsQv5247Q2s10Cu3m
T203RX1edqKwadBiNzEmDnjCnkFouRAPEgqvJFV+qgnU0dACsbZzdLpbhBFX5kVu
ZaGOmu7jG4DbDZfgZvshwlQwiptAq0ZRxBEgOvoJ+9thfQPQMJYSxkIc7kCJOIcp
+tgXfCFHAvE0OGSKOTrJBvi3N+jkQJK1xlkmeNYyb/DYN76x31avntxSKURnWwme
V1MrsfPU5a7A7l9MKZNUf/y/bfluCWNOUB/2EwnysnFOe7cAKlmDwBFlZsX9Rl3x
Mw6gDREeCVB6gC1M3xRpho2EpxP0QSGTe4QaBeGUfZ0VlFpCQCLBdBoe980EkDa4
khfPxii+lixCRGoPwkuYMFdQD9h26RCUTElxPazl50K9B/EM8Tym9RUtPH9On6G4
6R6rakj36WiHlxxwFAZ49R50WGKBiV4HR0Ckc8L317W8xukB+re2jD/u8xsmfP2K
8Z0gQK/iSVZ8UFJPfGjeHjhGe8mnZr9htCi8XZAVwmTFDNBGk/IKBkUc3QhPBx76
eAG7iM2Bw8mNuWOVDIteIxEy55pNfJkJfRG16jiLzuQle5w43nX7Zkn6+UZ6GQCQ
tCug/LLr3tKSXFyDs/U4jjAw8gepT/NetiDt6MRM+EDA2XLIHU8EJRaEz+JCB1Kk
1o18kDNfhM2YpCMcDtQ/HiNEGjnrLp8z78QMMZ3qubgxILlAkJj8lwPW2aHwpdJG
wdKfjKpezdG4ihsvryi7SKIdCvhiewgTcsrNjEMMwZzzKBpf1/oVVhzBJVPNKZcL
YX5n1yIZZ4T0VGGFoQgInRmctj9meDGk/B2EhDphOI6w+6Xu54bHpNEAQPCjrz21
6+rXk9LVD4lIxcejoobH+orgniK+zl7gDmoRGfDoOo2wvp4g1S8/a9toIVetEte3
6oZQdcMAhVltmx8N3NyeCiBHfdWFzo27qiL9hVDB/OpTxSYjG0G137o2P8InZVX6
DCyMv62h3Cs51BdmRzH/Nmts9Ipetcb+W3alAZDGf4XWGGN4IOgzdJqdzYxSgKgJ
YxRidMQbW5FiqahWejcmLMoF5G6UHx3qe/6Jtf1c9Vtn2w/4LiZ79ya8t+By3LyU
l+kIdJ2+/0KrQCW5x/6GEIUXOu/rSJR0P8dmkQSTuR5ho6LuzCDYV2511pi2u6sZ
TOW/xzJfJGidbj7mlaHM2q8sDlHDHIDiu1tz7cblpdBsI15Mi0oGITxBh1BHTTu3
pu8dxmyXjMY1qQymQXU3kObfAzMdxr+45/dSgYDVkEBJ8TleNJzWZiuaNF+K4n4z
VIUTX46i8/rk19UW7IeDaSZgoFJix/x2cXrWjXFPaoiUD3Wf3XMtycndHM4ccMiq
5dCNXFpJf362IcCoSXNQdSW1teU3tSywqo/y+FUkV7fsqIJIRhvj5zTc8xnmpYP6
KvS1zUxs9sDnnKS8amlJYf/PoRVFOTBv2vdfznk923JAFfWQGpkyIlh3LYB8ocN8
uh95HolKokXwy3OugW3BA7zg6kxfkNGCKUdMNYW1pmsWX7PVkFujAldk/s/D8K+d
4wIDF01eLLu2O5B/sp7U9+6sXGcPBi7OJkP4xT44sPaYBy3yB7Igaj13mHm96Orz
QsJAwmr7/QrgRkSLftDJS/PuO1YA9B5OCFQNL4LbNncmsMJP10zgbJqBkG1Xxrvo
bTyizEPAR0nSDAiyqHpOSNFilVOtCqO616bwIYX0kC+ltF1RvPBepf/QRVq6cx08
qqEH70ZpFd9OS50KaJ21gtydUyLYKgbrZBHd2rdWTRjuUBfwtpy85Y5PPUxvE2rR
crPYTZ10v+5QDJEvlmxqPWwNbP/4il2ms5HN+jKU4yAId/K4b0uRABeYmRv5qivx
ebLzfJPLXqpHlJYLH7qfuK8p3nnhp4u6Xf7dmqDhd1VZGjfUkXfWBYitwaO48jDH
8xNcB2cUHsaGz3pei2nLSXsxcBKe4kQuUCl44dupGFURzZGEX40Vwi0c0RqwB247
naUf+rT1dXFbCVRJxXK5iUPrDhqCEeLzsFQ59bbh9DG0VIYUpIcmrClPoyCB8oHL
bwcivmIbXPvqHsxwh3fEqzG3EWtNYZRQsKJFll0KnEgdS/3gvQuE9ToaaGa0ksEX
b0Mdb5p+OnTOcryZnTbnb8BsW4D2fPj8ex6fWgu3AER0tx1YRqNAF33r87VBnE54
SW8rcGuJAsMcDLGQEtNircpvxLUr7Xm3NEZQR15IhBYRkASHdkSO6GEAh1fI2hxJ
OlXqBHkGv69wtAVIdgtE3J0tEnnveakIdx0tKQs9830JwHYj095n/6KufMrS9kzH
sWdKFRTHyNi2ZOzIvRdLn4fuxVCQrBr0eiGxGwzAJXFfkwYivLiXgfhEvADaBkqI
fSv9XxwToZyehHpF+qqL9MSaRQVI5CbfrjbVpeS7L7IrBg5q8xoTyvMwD0JKtxy/
3pcxAAAT7IHBtdLLnp8A9aiecFZzI6zwVazgV+xJvi7lXnfUXUVBwmoZmdfrDld9
CuWqGKJWLwdm4YfVCBJT4oBFP7iEehxgWMaeWsR9vLmtTdujd2BKR1nS9cLFjmEO
DVyTYMxYlZfb0dLmel3aTLdxYvNgENnYwQUuFQ1Z83S6Scl0fSAufCDJWJsQ3Ub0
7vgexBVSXpugngoQuRyDlZJs547A4AIu0Ccq6j7ZKdzkrqWhQTeqJWRDYd4Js/jW
mUTiRduoekOjlOrEkVEoKwJuT7ZmTftAHWATZUXyLThObMliTyIMFANYJFQmzsFk
X2nNdgCPPe/3rNEIlwcK6L3GeNU8HIv1JvNbpXpoyPvtgY+tprSjzWDgS5qXIYby
sZyD7cIcQDRkw9vnCPGsc3h0U3e+W8KM00o58sYk9y6J+780J7UW2Z7XAO+k5ATl
LttjegoV/9PS1rTsLguhml2ceQRYT1WZNUkpZCtyqk8NLx4/t2BJFM2sRPRWvrYL
BhwLMT0Gfd5zEgZPsmq4N4r6jqioEe++K5lo9Zfq+3hGER7LbV1oVyjsepnz9nWB
YxdFY12BHbQiQoDG1/Xyy/w9Q6GLX9e+C1WD48v+GWYhwlE/F9uJzIiNWonudLHj
WROxut4vOqdAEJks5HxoqTeyXPBlIkesiKHLnaSRgFWxEYG7VgbO2mqRb5DkfDGr
FzcdwGCLgknemMlfCrexcoK4PuTsAX5Ey6uJ1E2L0PurwC1GPa2pAKv3IRaShbxj
hqxWQA9KyZzZTK6EDcbiSqudGeKFq911tWE1VdYX9r5OAfJaWwIRsP+5wWSvHmmc
JqnmWn2cf0BHBlhnovummQq11hsqvIlOC3yiQSivEQrgfeJGpvjXbLHYcYpocsjb
3vvBSZv8KfCmP0XwEu2HmdeGykFBGkYJiYkF/cMc6ST0PBk2305M//THCMqF/FIP
XxWQlRVF/nvbLHv9qNgdZ2/M7OVoxIbSU2K2RreMQRLR//8tfmsVMd/UCM9DG7XN
RQmugw03+Nu7Anvoa9hfgaACqXYYU7syZbhwDv0qW00jsVYNleBHAXz3YrmQg0qP
9s9NWkHyKir4YGuL7SGE037vNEQO2qBWw9X4Yw/6brcP/aKSbjT9O2OM01HNCNPM
78QU2xYw7j+kQQt09rZgkYktrwwCKZmYf5azCY2mLycpUV0xgfS5alO+9gQnpWH0
LwFqgH6Rwx33BeP6iN81KSTJvB4uqyxSx/pQhJ213w9HAlfOjJg4Ph+ocgRMwqAn
MJSuatjBv29w5tSYVMCFMZdaMJLtf7ok3N/zOl8uRi7J+zlolSvFnIcdvK5ghWDH
PtCdo7K/elA3QrQFTLiR5turzU4RJrhAX3BjPHWQwFPP5Xt08QQMu4EMEGka5kCD
8RTQF7VthtYxaLm77mEdQiZfLyvQXtm//eDcPJf43rQCruQ9xtY91K61FlvkemCd
WkLC17oQj1/8SScBH8d0gjPSDo/5xk9hHpH9VvzxpT2xi0V2WDls95jXLGVr6580
z5uWHFd8JKbkkl01pydkylDEv5gyljkX//FzZQucMbxEiZRmO8C3QhLvwBE+VfR8
AqgBttQ4ore/8BHbXWsBzTUz7z1wTclQJepOMe21ENYTmzjtQvhCWDQrCPbVFHwQ
CVQUbt+v+jhu6sBNyTvHDV7/VRUFsBiCcr2tgQ8t4ShhOsBv0ELuj+Mf3LyXbW4j
xlJQg+duTd3Dowi6sqXb1I9Fw2baoTlPNwec1jgQ6yfQr5m5VfYmnJ9h1OkS6NVE
rfQCHpxcyzmluitU4QO4ttY/xVb0yNX+nem5jFT1KBNXK1TdjV/84ypKrkLU1k/o
QJuxdBVUtYiJKojQMYOjI7ZR6sYzfqkSA6PDMmXMJwc8rklt3VbG+LNO/ZuL+oO0
BnMJw5bDGGtVw4ttrbqBpLfEgC7DNDDU+YseE0AsyEVmC+yQuIehbXLX5+sgGckV
AUAedIMorX1CC7We/jWFkJHoueXV32snmeLWpbs7X6RuEVeR472VjoC3QgknLKdk
LRGwVfciJAgSj77oV5rhhaH1+6gps1jxX2A2Acyqkfy0nrLI0sbSEX3U/9+U6HT3
JqNgWI2dCDYWwZp5m12coPwwr4HWYkKu8BK8+rgihL0xykoh7z6ZU64eYypUwvE+
JcT1+MXr4bS3kRKTdL1DoB0bXPS8LMBUX2bGu9p8YAuH/oB0ezqp4TG43sjOrKIP
b78hPgak5kMmt4RpP/C7JwDYOEPnkpPIhUsMUzWQk1N5i4UIE7On1vnMUKC/zbB6
w7ajZntiZPQZFz+jJYHWela8TNeBsbtDjGggJS1wE1wPQHKW+j6IdDX1yJIo+Uaj
3Lcm7L/oPAdgSv68eXy544VNny7btFq0WGjzuVbwOhYmeHQMwyzjXwu6qkiq1AFU
Pp2zkiQ+sS5tqu1eab7/Tbe6zUubbRcpIoERFxG+F8OYoNpKZbZecRYPVyEg2NSA
L+dnx6Xx6S6t6KIZfK+vkqKf8fH1vXGU05ufF2GDDVFAublQPXhM8KzAsEO4z2ND
8Jq7ZJHBt06YJRPJRAzkw+eguMxn5OPSakaE8n0ETkoFfpXwaG6N3B/N7sjo789k
TSdsbpd5XUMaumo0QY6PkcpDBL7Tm3y7dRuif9BgbkgLX7W0CYZkoLEl6J8E43sc
mBMu00nV0098yHIpTiFLJ1DwdD51MZSnErkL+c+9bhGYwsH7IjOeIkAN1u3crdhq
uWYcuCweiGrDAyXdFQhfrLgJsskEzHWROs/74SGlT5CMXmlS7J/u/1Stt7FYj1VA
vSvhbeKBRnXvOXxQrsJvmKjmZGQGWQTVcYmYfPseg8lc3whH3OT56X0JxGBCy/Qk
klaqltzl1Bc4en7iTXyZmE5Xi2v96M/nlDOVVSxlIc13sEXkHDCzDCznk82HuqzS
iCW4qtQUsP1ySyoIvxWmZBD/yaSQ6Dam6xk7OpDtDengBfxYMLXVmaFcVa7W4OQz
lJAAXdfQe/27gSJpQvXYXvW/Mi5AENgsn5Xy16DnNuXs2DxJCDcLg8sCw/ZLUlzJ
qFE+4uPhmFDDKlj37YZofw3A5Wmi5RgS8gI3fQ3BbyWHOHAcNzI7mnr5d5uSLLo1
wUA4LTMB/J2WIhM6DDNOw+j2J/WoAG3vHbbFXXZ404zUPrQBNJ3qQ7IN8wLvSeVg
mrP8u01Mr/2SiNvULsHL9S1FCEXGGyRaa+AqBQKP7QogMJVZvPiTLPjjOy/1Mz7I
bKKe6nTnFrYTRKnxJQiQTEb30LKQiTGpes9CHrzgygEuVMU6vn+DAufkMxP6YYfK
Kmdzm6RhQ5ziO8WHysCE0Xnu6BR4vBPVGfI7MJv7n+RjPuDuS1vYvftpJyoMxDVd
PFtdw3A5yyuLRuzAv/8AkeN8h8PuUC3IVWRywmMerW/ME5lIcLeP/30iNkCslU5Z
bO2qFhZMEPFmvV4MNlSGFS8SQCKvI3HOufRtNxL1oWumWBkbhbqDXbiJ1sEL4Vnv
X5juG3/Vwa/X8qf5lv+XP6oSdMSkJVlCPUfSsdvn+AJqqh7u6ArX7PGP4uTcRRU2
Zbjq2FtKXAIJjheXGwYTPcM1WPvLpLznt/wt6aILqL4bKhGINYKKMtaT9FR7tmUN
m5duufMo/EJHcaZdMRC+uzK9cerzctXTR50B+ut+VMjuGyetMBP0BYTOSPi9IbTU
Zs4F+wpNcd+uaIRSF3oyYRO9Umep5O1FMWro71p6brXXF/uDXJVfjp8Qwzy52Mp/
56uroNK1sZG8OhDxkI33pIrjJwFOyi8vlyjIUeQpoUx3fUV+559AyJ5hy8LHgsRz
pQTdj3cAr8cDTMF8z4o2Yy2G34QzFu/NGlnk4VgzyxO3p6HIwoN+qhBtjJkmCOaM
bisZzmZLOfLkcUw8NpHS8ZLrow3wPI77+8dQ8B8gAgkTMLcVaRlpYzFklDO0q7Po
LdEdoc2vIb/akHQexX+4IjY+NgnqOCsmWr7QC2Ma8f8Snj/LMQNGeDkXwF3kBgZ5
bCl6DTl3BigOX2i9tKYkcdKusza2VNzOn0mWYYM3JdJTmBB5ymdGi+8NftgItwUe
Vnalw8XqZzONTZB2DjtKXtzi/TNfri0FttgGQhERNv6tPukXNpf69kHDQcJFoLl+
5GQYi2PRCSMwBk+Kxhb42Coy/pCVqVcWRJ56xy8lb6h5C/0YhtRWvG+w+l7SGQJj
q1KjkRoUPh1s0IpsfO8vuv7pFr1p9YTbfekpdZAaMWZTS2S1e68DaFSrnuC2/+UL
UFUicyiR7Bi/rQIncTP+zk6NKz3ely6i7xRxSGFm7z+IZ92UdrCNqQVa4q1SRUJG
46wIbIg/AFG7yA7i8IwvHv2vV3d+V6shHLRcg+maHNpvlRYJzdHilJ2g2Up9Gu1q
GF6rFX1uj5DN5D3ZcfuJ3SI5yfrWw0kr8bXy4ciaQlAqOlGDmRJ0dY0EYMwSZtoA
lLUH8uzB4L46eiYUKB0/rzlHENr1fB9XvTR6gabyxrzp3KO+CnJ2aQzWlF/zblaX
z1JH43Wo5GoUWfkturI5ShKOgo9OXXEcrPZJuW8PB0CK1C9fzl4scgKIMcbBVgVo
snfRx2xHO0pZcQ5a9pZ3fKoaR5W1O3vB135ZfEeIgE69j5oaGcTLgKa6GTk0fCSS
tJj6YmmJkQc3bbe6FOhYIqEMFpKuM/yfbgy5nz9uMcFdItJdgPs7IEQZl1LX/Xyo
xoXEaaIe5b4fFBmZAVMsTu+cOZ0Z07A1g/jS1Tl8Zatni6me2HfluuWjX9+ERyUE
RA7T7llYEEqGFTD0GS1biUn6VQVyPb0SMVA3UpwJQmnvrWaqTkrQs2G6BMcspe+q
kpwO75TqarFbQgmJ+5zTugsCubqlE/e2iWBcJ+3CGQ6WSTrqQ4k8lIj4Zs6CyTUx
wS4y7sK9kr0xGYGf7RQ6jVjQ32YtoZydv8x8mhDQygpSs0HNzi3WlmND2jLZ2gNX
b6PW48/e6NP9ptLfrmgnqAsiXej0U+nRSHi15HuLcyrpYYf0+r83/u/X4YiFvn4w
9eS4LlklOq0BnQffxCLpXaWPB2IMrdkIeXwWDdQe1mhDVhV/2XemaG50ff8O/tJ8
yizNAzinmcAsCTwkfwn3I5YsmCf4JecsET9Yo+2ljfIRHbLc7/jnrY7sbe8KSNfz
ItF7ufBqxXdMqLNpy/VtfJjQniy5FL3C341zfnAKqk7SLVcO+JVyhjcRHOaDClsw
aLzxlvMHYX9PM+Evy5NxvEqKbMIdGvFkUl1taHvyq6j3f81NDAkC/VglU9zCx9tS
sjJkEZe0S2U3iYAs7WhL/I+2lTvP3TkFvG+XsmTl/Y0tpyi3I23ORAY68UU5i+RT
+CAvsHZpzJ97bnA6PEMFOS1USHR6XuBqfAUYtUYl89nFj6qmwSSCNMfKGYSA3eYW
tNncORKERLZsEPDi+hH8LuyHfF7kjwA3zs8rJjS5+RmgtY4ZDPzDx4fnYeABPqWn
6nrtX3WR0N0cOdkrTRDswyXUk3VSN4qd7+xyfOrSGlJM1gDKzpJH7PWhG6xidNUZ
u1e4A2+LDlSlat+I7i5qlhOMi9giESSy7aGvHDlSrsD2oe5pbvlN20UCsMmDqU+X
F8rA7RMpVaIEsDV774R5GYv/a8VdPuRD/hlTntuoMfFxNewvZhk6qI8FUmuQkaAQ
0doG4u5yZWSUGvorHu8oGN3jjXCTluz4rMhX2fGD3R4/1cQVOWyYraO9VFL0xjAm
7RNAiz14dpfnEvI1Ck3ht4urBt8gE+luOdi1kjRfO+LPhLXELVk+eK+Zpx33X2BL
hjYHqtSf3sc37IU4lNbxoOGKXRWFtbpduzfpFFLzryKUQtFhkRHuQRCtHmq0tcvH
rtg/6Yy893FLabxSQVlPdr3mxAkd6LsLtaGc3iURQLu5wlOpI+l5FMaZHDeO9WB5
UMSAQWi5rILlXX7OJ9T5+8/XN4t9HZST01fS3/cfxV8NjIHo00xbW5tmAuQReFHP
bpKxeE5pY88TU1u8VG8FduL3vBNgYxRt0I54/FVjY03xZ14m6KgmbRB4iwoPqOcq
vTxazTPYytrTDgSRYK8GU10jA+PLc8JkUR+1WxpxTVjKiI6zkRuxAePTfCIsAYkw
ySAZb6kK3VVLjeOBIyvbVF0wtmYKHVnzGypWgHldTm7QJZ/VRwZciQASKMVp5/FJ
D27gX7x1QcKX+DDKOHY7N7JY4CTjots0mO8pUfwtiQhOsxeEoanjqkv8Az9I7x4q
+NqmQL8lBxruXdMRIVczWoI9VcRQ3TA2+daF/PJpMpiTj/zl5ExlR+RXRFBw47/y
11MZ073HpN3EirJVH3wVQNqR3pZ+e/ecf8n3rEwQiMQDd4jkPvpnPyd2saoMWqYj
xOaYmdRCspDWKtPn8nqgnzxJltaa3ibfsqDqCki1DD6mZ8eMSgUkwVVd7sJ2wu7M
V5wWulOpA8mPuNNXVR5t06nYkchjZIVJ0vmUBIFrBcC4YYUdUoA2sr1e3KyHGJ1s
vebh7V3HlZkwxaytprGcthrZqmp0fppYgGfrh/dsRnYWwdcGT3yyqehxQTpHYQvo
OGQRc/L28QAByKnlUDBV4Nm5a5djRslW9KF2CUYUbTvYwVx5UZBr22TH8hqr6kxW
m/HFBOL6SaNkV86hbTWoPt6dO6BWiAzqUoStI5hEDvP33rpYrvbiQ3Dkk3z3VVAq
8pekEIULaO57ZwIg/qzTpkOiIQCNACeXAOOwACBERRtLczbtBtTelEocMuHYSTtd
3QWuUTkdYHPon9ptZJJ8lztnGSTUYmTjBU1ZPJrnHWdIEKTgxKrmRaRMwWDqU0Or
mwhFBv1CdFTrMAs4HtSkmu95YS01U7GVv8/TxbV9bmy+wl3DWOYKI2+WZ2U+SyYO
/lQW/N7CXwg2uWjX1fmuBd0CHAmpolmGPgYJau4AE77PaWth0+eU4aLn8gjVqlho
jEAUEcSWV79N4+xSY6VREQru3hfO06ZCcpQndKcPtbIQ7CfBfj1cjqqso7mpHAoy
lrRKcwPcvakaVWUdC2zVC64yaGXCFepC0PFrJwP0YxNM1YuLITzsQCF5a86snPIT
CNLONwcR48Vinx4mvq6x7WaJ3ailPt/m2kK5QAwor/uw9Iqy5zcRgqvvkK5FHpA7
Kqzxfo+VF+IL8P7NAjxxOg2Xp9+N3bdCBhBJdFuukyyyqmqhMllpeNzchtrHszQ6
nLvY1J4ZhwXyT6qHw/cl4QXK64DT60EcEmBlc1GINHuXu5UEpXqEHETwcJH+VVXg
7/nk8XU+IqSDineaEaX8uGhyjMB9zhhOB3VCE2nMkjRI4rBbwRMnm+Hf/bTEq3Yh
IBKQ/eUZkUx4zPKfCCBbHwWadvIqsxQQxiIsg4bRmfrF5TzS0vVMd3C5MHp0/CAw
UVvkkbwcZalpecUeD4k/jnLABfozMioUszafQJ+NlMAASN5XvUuQczQcwtRrM8U4
e7EmrLV7Hq3VyibMXGRDhOirF0AjHPdDUpxYMt6ZrfV9eg8F7lVlLVaSsQXsoAbL
YYat790su5aeZGRBr/EzbLb/doJucsxIlWTYp48p26TfeQgN35QUX1t4BQLMMJqP
rGzMgMAfPl9Q6rKY8n4uRcipiENTMwbAOd4is5NC60hrR3JAcv9ykIX1zf+Mgo+A
1oQ92dvGGVD+/nIbNOxsc0W17hvoEY5YO4WQeuuaP7m3aAguTN+4rJorcrCTxeNS
lsNqb3HvIOFspcc2THLn/0ijlZJLCuAUp25i4Mn2WsOSKSv8vU1wLMaCEEHioZ4+
3Z1VSz5vuN6A0n6exCXpY8+JpFmAi0ZeIFkDIN3KG2uLYlAMm7lUeZS30ibRJels
DWr9zT7AEEHC4zVY4d5RYBtt9QeaKYpGrU8idcfulSHnNDjcEMvmU3RgWQ2xxI4W
8hd9RQYXsM6LIc/JebHfibDQADlcTvADOCZxikKjoETx5PB07GWP0L6o3wV6tdAo
1cpWroMoqKE5d11JIzrhEinCqqmh3h++bygUiL2vm5l0L02f4kOeHiyO6yifVO2Z
/XAKt/i0JW9O7dVSE82ETUF5sfzi1MKnJ6hviCXv0RsC5hIFhXry0GzRqiBrJNl9
rufeY5gU5ZqFqBERhDO7nD5YtDJ/oaAppiGDgsGpUxjB+xy0XdlXiktgWaGk9EtG
fb9T+RDnfg1zS6K+ltvEbDC4ohxH2DieINvts1QEtOIn/RqfURLbeoNuDC2kTchL
RCKqMdGFQgjQdFbcttbUUHbYwXtBDzHQMONocDAFZtt4KNrOA+LgtNjUveVXidGK
zPBKqxphFDqyRsVvpsMvCeJFMn6gHv4SoRTQZR0+lFExO0bDADKJW678OybHeOxV
5JaP8LxIxYBq5kaYEw1UOmVVLNuxXD5Lm4JdSEGAzeJbjpTs795FT1rrVAyn4ET9
m6OCmgzaVfXOTeYhvraw6B1mVycAhyte0CneN5mGMkhfOQvBNpPkBHuAppfxXZXS
ObyN13ShFj734KA32Si0IRKHx39IZYTZeIptPBDo1aK6rRkhTZzjtLRUfqG6IJhu
0j74PQaxa9tTBtZjpbnunEIBc1O3rVx8CjDGbQ3m2cctKDYMfD0khPQb5ZELxZRT
IJOZAM/gWsNOLts9Aym0wTEP9HFtQAtD2nt2U023iRh2FjiOg93iEtz6vDG+5Vmj
zhOzPMlf7EK4Mj8WSC/hs660w9a3jSLlNM4CbVwIdUB371Cfg8ITJwsTdnU+1M6v
fh2sEsvNqEEFepgNdHrf0ANZj47EILSCgpp53/W6bOxWMEp0vs4UT0nRoF9Qk2zO
561Q3z+mzvMJZiMOAzkOuDhfGTYf2xJUL0ojZj61PZrcs47bYtt5Nxs0+H3UnLyw
SF+Vu3D/nTNUs2NaG5d8nZmQnzVOAhDpPnXFDASEK4faQ4x+rFNhNt9EmvmYYBkz
T8Y/q+3qtE7FS7NoRkHtnY7TNwp5/QWIjr7wo0sq0foH/T9jBhUdLLqzDpjA2ToD
52W9GMRVttVBFeYxJt+ZmshV6Kauxs+6xCo1pHCdXmcbEN6ukinNQXvCZHBNdu/H
t/b1mahU9CTJ93HLgbZxrFcKks21ePfA2jiXq3jPp9GS9tLGfckLdWBWNpblTWre
pSk5K6ImQkduH729MsQBUr6x/BK6/QNJgTvyO235vXDF8cUIMlnMmUqEZbF11QhT
kusanO+0SQgYqiMPQv8q2S7XPU4Z6px5rF0PRqiBcpKoeWOIMNP5CTTKR889Vij8
Q0sDcuVcH2FgsrhomMrgRHJd9Ba4YJV5f+aERRKToW2NFvwnlP7yKjS8qdyoPy+6
Ho9eZOkx+ZoGn3lTJNhqBwgODy9rvJ06LW9Xjk9iVl4l8Wc1vWqBT2/H9yBhtJVQ
ed8MEKVbejEMsecOkiz42vLGQzc2pz6/DS2BIRmg+Lz2B/3S13ncSzx3smDBOstr
xpPc5BNYLkGUeNS2KeoxkSsByMageLHZxJ7ds1IGck747es3bxwwRzZGBg2ZIFPJ
tQ2MhpKPXsOhhJ9Z0Bnw+QatMnF6ED7iEwdzR2KMbT3GGX8LNkis0rf6HZyHab85
O6QVfNQYL/1FfbasQqdRab22EG80W9S5D/4VNKS6dj/C9+kyrTZfVo+8usrEA71Z
uzApUaazwfe4/1pSB2wYBpyUBfrZFsMJXAhYJKBaE4MhzFQfrYXjsCjVRMj2A0g0
qC+J5ANRU87h8DkxwBYInqwnNKgAVsv3PEQ5AcJ/2RlKHqmCVeeJ+b0dJmEZczH8
dvz+flGEJkjCwR6pihn5wRA8ZFgizLFFrfM2YlEjWN6kpeopJTMW90EAzuP6hIRN
J4OHBdk8HKIyegGbx7qce03DCPu9sKD7OxOemL5g4PG9SAmK/RMo5ADccU+sEUTU
LbilhrwKg0rgtixYAfCHIgBQtsA9fychJTZIh5uIOGXxHp80nBrAWikyuTlTII9a
UO/c8HhVRTOfpQMVip2zFMFPTy/7BK7tuZrZqjMtshZh1Isrj/7UeOx6bo6RKlLf
2HPzdgjFsCp1HAl5fIsMPyEN8UUW5PbPzoC8ubgG5J7JV797oWfJ3Inq4vclqKJn
LBZfvn5GAClGslkDutgBNxwDf7unFMUfbCU2pZWeI2Gka+9pwTIFw966qIyUIftp
YsHqho8w0ACSpGT9s5J2CoBb3mtrCFkIvNKakyVimbEZb6aaJfwCcveB4ja8vAta
Y0/Re8vFrRQ1ohO4LIqilMq0BE1Hep+CbvAG/YJMtqWACLYSiqr0evqbdAJHEPX3
2sKtwkI+I5u3Vvwf8ATECtzZ3leBYOAyu7CVwfmUWFUEDsXRK6M4YzjZTeJuPHdb
xQcDorv/24X06EwbSP4Ms0Q+DZx10Rb8rPwI5iVFM+DjjBs+AFTLxypxYBe5SNvF
ACWNhrG1xVu117TpwZHlDv/Ax4yXyoaWy6ehS5/5I0f270NMnTNXQDOuqeEzr+tA
bysjYjW6/SU83837ext18zete6w+u7L5vwBXGNE9SIpmrKqcu6pgy9zk1X0gsG5C
RBFch+zGtkj/b+9hmKTIB8zY56RYMAu7UbhVhlwbbLMfXlGF87w/4UXPNHgIv3KD
CQMd5wL5WrIVyqCKbhGqsh+XwlPpPCTzxy50cro4lpyQrsithBqtPpoxj3QuHUGJ
0suGtwiQdASB2CPn+nQ9AlY5W9lyS8pVCfmhb7cEHKLaB3plthtmh0pGIFO14OgT
YhdFcagA2b5GB9IUafmZ53nJmYI2sGdEF6AcFCpCzQ3nFmyP1knAJ4HOuMXzm54E
L4ybHo4FVG9kvurQYN9Fk+H12aAnh5f2f/78hQllr0gNHgMQqzFi1tCYvMg3DiCi
9/p8IzaLIet5Gk2dqgE4eAz1Kpz3NbvwoBBw8Ury2Z+p01PzLrn9hGZLb4jDw+fp
qQ8Q9EcoseP78zQHoU0001/N/cASvFB1mYTmhNXCKwzplBDJQYo2dWeZRtLP5/4Z
DDmsNZYYbJ+mdza/wYo0Td46aUwS+su2xQIa8/44JiyCMU6jQTDwKrHcZ932UdV9
dypW9uK6meRmM/dKwI943rh/lAzBLQsEFdaY4ZLZ7mwr7IGzwAqLJOcR4TMPPRxA
nki7d0O8tDaAixBdL4kXgX1AIkeO0jTVOUKsqrMfchKfaab2N6XpHK3GnIcslaip
ZyFNd28hhr7O/YqMmYxU8xgbkQQO9+dHjq3OpF4jnfeRVjuaaksZZrjrQ1NyYoju
Q0f79tJqVe13evxdEuLK6KyrJBQNyvEZFPl3f6pXIJuiBCALMMC79Wc0oTJ8HfQ7
HrGCt6lFe3jQfKSMiO52w9s4PqQCeDoZeQQ+bO6RIEqV4MwpBaTB7e8zn21gPQTJ
b+ZLxh0ljcc49pUHXSuFMhdwPMeOB88MB7v/aAQOEKOHGT/7d1mV9/ssGJ5Zf71S
d/bNWFAPTmL44UmY8sJpAnoT7bt4QrM3jX4UwAcvWTr8Sk/+Qlw9U3HQ8IdmZySs
AU0VCJf5dD4mO+N/pDZuewmPhXLHHLLrvbYYoJthvO7siYP6YMWMH5zsLvKLT0vj
dFkD0JPCOBwq4LDjxPWkrqJZnA4jvOKhRDwKASA7OzYBe9V806FMRFXI8WXE1bq2
vlO4Id1bJCw58EjXcqTUSwZ47UHdB7vVy/TIz7G1DjOl+ywP/WBVX9YLt76RIN83
BZ6JN7pU9YvaQHhCSpnhIxAbQ3eD89Rr9CP05ZC9jlu2IjdXbEq7TS8ncO4uDL54
u6XiSHk/cvAEQaerXJCiaGpIH2jJpDPhsprkKNjcvZN37nRbszJ20+VEqevcKa3A
VN0nH9JUgiuXkttrhExPhuu6M8gFSJnA5nxKFWCYa1IMiUF8TBLdw3fYm9xuW9tq
b6o/QtTl+y31gYse6Ta3bSm6lMK16A+3G1HNvNB19us0HWdh1D28HhDbKh9k7HDo
8kcLQis2hTDFHMKJJwX83I0DR4iafsRzZ7TfoIgLQG1a3rEfmwvhCPMIY9P1VK8E
vA4lGl8PZHvwBmuo7exN0sjeGvwpSmc8EuUO8tRCUt1E03PrEsru2JExgurmDlKk
/UaHby5HR1YxyTNcbH482iKNYrnnOynKGaZe4yqpysB9S+6TPRC0hJXVMlumrZzj
AouOBj7hDKou8dHeDK81ZsAz4E+G3lPELg0JtMitOnX0rp8xnWibZWejiADlUgY8
hDTpQ5TPxaNigEsozocaXD9ngMiIX1opVxb5R3jirynLdcjz5Q7aSGEUu9v6JefR
BJgS4xaoxBB8y0SCFqT32yNVNxirp/Pq5RQza2gGVVGqMVxDZBXJa0PoNGIGhv1l
P57dMwsxD97g+stbfWxtbv/mehjsdo+0uLqcKVWnRBbMntwRTu4XtmfHJBCNaJrR
clUVZP5pWE0qGYgvbvLV5irrTEwPiRChw60jmlWgIZNVaWXW5/AAjCf7g4IQab9s
Yr7agWG9gEZ8HuQcpizELPL+nkCpGPzVBOPQ9FAyPTep35naj35Th3n1+7DBzOJs
NUR6SHsXEwI0oh9dfoPZuV06z4E/s9TzOarQFK4/iSAJm20TdA5DyEzU1Ie2bseE
IAHuGoRhusJF0R9i0zdQic9UOUiuYMNn7jTVFJYgF4B6+58WG45I5YmFfZUyTvi5
q4KFrkKXvL9o+zcprTupN9hxtl0qYf4uFh41CZN3yK19hEvjKEG9C9ME0HWJvqW8
mkuogfleXm633jgoCDK5eSHKMW2+xu5BDQjeaI/oTzxiFdLpHGGb+oiKsk8gnrgb
cUbJxrpVckJqauK5j4CetHOWQshSZiawzGOWEv9ZiMMIWfwlVijGQbD/kru7n1Yi
TS4KqnDCQBKD6zYV3+1llB7e025vYKj6+CLAx9B8E0Ez9iYcQUa+bfEgqO5Hwm/y
S0g729tO5JMIG9rq7GHE8NIgW91W/6GTcVPZn0wYO9IO0wlq2Nh2ya6bnCokQbcS
IeG63994mKU7pqaRiz1MFfO8q4njOljozENLbaRKreeyv/Ev1ieBe5NcKfgxJ46P
qgrFNi/wqqS0YQ5PoPot+satfK/AjxiQztDcMLNl6qoYFTkQgp599/7iN5l8gTix
RkxopRWUtdDqG91eBjeGKfqLwvdP0rrePnUON1Tss/6Sh8kYVpkVr99tbYySogyU
jmfqrPbj2zhocYLaxEqgcf0vPtV9JhX7Zoe9aBwpxy8Tk2I8MWy+57f6lhZfI6Dr
ZU9kOZH4ZlOj9kTlCZt7CKlcOyy+lh4WvlcAruLk0H7S5kKN9mFNJRz5aQ04eIbN
kgrJTzFd/8JIEnqP+IP1wA78/4DXyzhULII6IAKnlsZ5P3iLGGUnyQ1NXUqs11Wm
T7ng4PU6ufA8Kio5vZ68GgtI9hPm0jZ5DRsUpNo1SJMU9XvGvab4/FtYtaV7eAUL
/++iHNlq8h+JCzWO2s8aE6+OVP59YngzQ5m4rfV19K2YCLSUsP8O5B2EIa1G084/
jvya4VBJZisYjmBMH/ifB6SJBvAa2Fg5QpEixYc/vf/BCvYTY/v2H3EJIdsfzysN
d+k34M9zZENiDqxegFnb10XwRizIAflFRxdMY1LwjlYc9nOL7ygoPDxBkaKWzGnd
ujvgyXR7KiB6+92+uwnvuI9DySgVkSyXscpbEptirTILfKdWkaId6xLMjFYwoGgI
qC/d1EfS7jFePVAaaAnHAwuu1H35/Mi4qCFGOx5W7b566XFHnQ8WU4ULuJn3JZef
ezxu9Lt8JL2chXQKI8Z1P1qXprDUtRgI6Th4z0FQy9yPpH7uumv0SfAhSBOIjZYy
e/tJtuwbs7scGbOI3rXB7F5oXE1pftXbJrv8am4G/sgeD5oQQNcn4sWyaTuFOKE9
uIiOfD6jTK7GYAgGaF1ANNQVx+K+YYgHQK9Hk7V2YHxCFq8YVN8F93O3OD9sR3DZ
mWLG6nVESHAoIHyzMkOzjh57p3N/gewHPPToM1vOx07/OGghEyvYkMt92k0H6nyJ
0zyyrlL0AXs0bXfqs00iffEACu9UntDpm39zDKCpGh+JMi2Ka+bKmNTGVP2e9msh
oHSs9f0qBU8bfb3Wle8XKbnAH71E354greHXKNacQ0239IX2VSBc0d1+eiTviceo
mm5cRkns37ffmctbmHYjdkYCE4IPHV2JkIFL+YeOsDSc3O9eozWjNRbhZzMAPcJt
RS4iBHzUy6+wkDZyxQz3pBtKPZ88uUBK6kbr2WapM6XpF20WD9GevaGRa/v/Y7Ov
jwEvB311CK5MfgRafOOYRNiBLuP99dXuJVbd8NihbZcpiW3iHDADYDR2wi98K98c
3RVfLWzMRLmSvTod6MptFS92BG1LZQvSYOwu8rWS6NO2hIv9wgZlOghGEB3Q9A9G
8gv1TOuS9NgGo7sXtnTRI+7s5mo22SHq5ABg14MrLpvKZ708l9a8sllzrb8ONdVu
bll2S2nYJ9GWPERMUEk5LFgNzLFCHvBBNXDEIX8P+zX7aKhapfn3rQAiymq7P8v0
AM1USUxiXRcXC+/seuBUa4Pgga/zPumwe6cATOo8Pl0cKWq58alFzIePMV2eyJjK
KJeP6pnbC6t9+rlap3/NACmxhSI6o2ePVPUjMI8vh4GDmw5vw2DRJxz9/Ws7WUPR
h1yIhRN6htX8lc4HZox9fdWfWmaS2IMY2dSB7CEW+5tWMXhxT7/ryffSi6WsWiCU
6RGpif3vC0yjvVQuQHu5fU2BLVMljHnKGmX8C5ZzRGmkn8UnQxL8lFCpYjo/tPC4
gP2H8FOw3iq5lefaQjkLTkmNag0/6YNYNILM7l9CdRVfFIDRJPtCinn2pva93TGK
wOteSl8e41z/aRQDTKMsPqcLvPH3BXUBn4nwIi+G8Bz3XNrTlgPZVpjU5o0xOfDr
3r3q9f30rDFunSDv9JpeuTwTXWno7pCsRx6m+dSKgROl40r+50+sJwQAFX1al90S
2N8wtWfmt8eiiFEOEVtB6YsdYXqg5/A+U3HUbNna3N9QTm9V+eWQzcnlrLPAem3L
0gyGKGECNUIcDF4h+IQ773Y0Gt6b6CrdX7Ey3EcUAIRY+0n8csfJA3RHgfYLDSQ4
5Ym1JPMwkZi9gGg7G9Uo9TStAPY3I90p93VmBjgEUZD9G/UTVgtiCI13+Lhl57Gu
ts3zscv+eQucyZy1F/2D8En2z0wbR0zjSPYe5+nFbLIFtJ9uILSmz7OuzAjgP7u/
yMvE/JLHAS/3LhQvymbiX32lVsN+6AbKRbr1n5t6AfK7g7jg5iaC/jxHjNEnmGX6
GQai8ru9EM9kfmdI2yE/Qg3EQvKNL1s+u6wrlDPl0ClYNZnT4/X+0Ex+WyfixDMT
DeIpl1vtIj5ocJPpAGF0ap9P6/wK0BCX0b0494OI4joh/iTlR02uV8UJbgxT1ntv
5XP79OLKKwVuFoT0QqdSg/VFGoVgzgVXJftQWx4r43MXEnI59DCHen2l7C5YrtkE
QOBovepBwXK67gHnGFVnrywmtdHqdXETA1LVfLy1vZOXMpwASRUCwJeSZ547NyW0
iPcy2h6dDYYMyL3HG50Tw8h5O/ziCROuTtGO3t+SU+ih5FZfngGh59D2AO8e1NUU
dyGJiishdktpxIvvMguDazmbA/zSUm3E64jzhPCYecpo1ZiwIOIcqpYV7SgWbMdX
rsUpb8LS/GSC7gCE3R6Yw10Zprk0Ml2c1RBX4Kf0ZomdQUryox+SLfHBRG5hLRyz
mppOf9YdFd8Z7+D/9257e8EZ2RAt478aVcaumvQ3lRvRDDoON9J5PzDzrFyjHKO6
Wrpx5ISe/JnAhVVXhaAWR0LB04qNWAHhyaAPtrczLkFXgHuLvEwSmkMjja8ikytO
GNlt9DrslVKxzooSNfgWursMnsrAs6d3plosMQ9OCPXaKriz1wwBniCVq0MashaR
FANcFmsOQV7X+Cru5Fkr+SIESuutdXjGdSpffucSAWEOCDSGFE0puDxq5BNdS13W
DoW1p3Q/4cO/2pAzYbyRXVVPNj4DOwXsBJ02KHMZBwPJ2bv66WlDIy6yY50AwGu4
A2evKroi3mUeBCD9bXlaS6HuRttA1oBdZ0dS9g7BX7NDBI1cAcmWR6BmxRixKCWR
i9hJLGnd9oV4rpI+jBPS/3LoZ3NWEoWoA4dxCDMaKZelDeo4bS4YWJW5mjbxZ4r0
EkhZQfpk7LbAWnYSut4InUz1XfHXs3LUYepqOPy//9y8WeQ7em9/vxsbpX3vqUTN
1sZ4N7ENJ/wlTE98nxTU79pzsPji1oPgD1CfcEEYKcoFn8+DnyaW026H6M4i4xRf
+/fbaPYHLLWpHf9rO95iYg9s3/Rp6h2AmocmH9rmdjKWmDrAmpdcDQLk37j5Pe9Q
MexBIZBIuI+/ny4e9jF2bks+0wQn3OyUj3TXywb0v9y8IncKwYcRXBOdkRBwsyg4
3z6CxqWVbIq9TUkEKYFov2vtZGhwqHoPNhm45ZilQkFr+RiDgTHEB1zHbLt37zZh
/XGNJ5JwETMaufM1SwCVqs3zepv4qemiGL+mHQe74WLjfejPWgy6FVjbcI/8om/Z
fKEhkpTO7++V650OmHpMVe8CC/oFcfL3JcOAQd5aRwNk4YjY/Bmt+43hbOFrQInF
iQxpPY+9LFa+SBQpHVBzevPpnKcrzLUUAG+gOGDW35H27LMf+qbQzB7e1VScCeoQ
7yGhX/VOIMBM0vyjaBABu87MBeLFOLVeXAtnpKCnZqBuEyZ/sEldi6Uee28Imgey
z6eB2CeXphrUwFU+e6P2EMeSS8KXxT2h3aKjSDFMxcTRyitQwiio9yDwXe3kipzi
AjETdZdk6UCGzEyfaMWVmLELKet7bgUalkXa8FuVjdsU60xMRt0LsEvRUOB+0uL3
C0+MLQkbP95KADXWDMNoE6ydohOjgAX5H6j/DmVXgBT1DI8VG+J7xcCgA3m27eAB
57qlkvMDAU8I6Di31ZZ35P7NeebD2VzR1wrPJcvDmYif1H39OH7lrYEf8Xk4iMl9
zSaNzyP8Y/A9vVnY18DQBMTQjA3sLtnM3UfLOoF8hwOV1aQ99tNTGdRGFgE4Tx9m
fAp2jD8V4hr8mKvRj6LqN/4PYTevTNVLdVukxDLlzLmjTfrJCdfJIegspeM+uRQY
nuGd6X/4Z2nkhg3SqDt5kbJlFR201G6kU0y1rypRYCCVCQnDwxkL7aLBNDuQdZmE
6hCCNgSrdOJ7S2A8Pv89/ykm32q5k9Tu3q06NVmRw/xF35ssSXYudNYlKU3j6KLs
I3D62AC2KCQdGYQKU2ls/o1yTF0F0xhyPtiVga2B16hDXBJkCwZ6PVf8NrQYCwAf
qk63pag0W8BtuSwSBl8haHrNrCbeZBH5wafH3prUA77j7xzF3HE2zBPfyjE9YP1Q
cXip2XD9w2EXDA8NPs30iyCsM702J2/9JW04MketSxoNNDx5nHjkNHth5QNDRjbt
5uPy69on195iD+u0Q0m3uQ0gDuo3qiB1BwmsMuD53ntmasRZKjcHXOFb+TyXhhPX
4csXoGw/C6vkUNXhG6tNjjSbuYqik/UNn84LoRrFbuuy8Jh0g0p2LooX0VPVyd6w
Fautcdk2tARqeach4mANJoSYVMH+QpF/IiRDWXHTSGmoxlJ8WSqQdiaO+Hd7gdI/
YhRERCuMUXGajr5efTn+MDviveziPq3Cp+cboTwezkxr83SblSAtUh5k+KhtEeZr
/X5y2I+OG5QEd9jSNUD7KAnlZKfsHT8jAYXzCSa/XEfYQTtcht0izW1lEY3LqvIY
N16ZqVG2qkGK6AvEHi55cGq9xv6TdHG+EL9f6S8kamvHM6fdS6Dh2ge1KoCvxfKV
dzLLV3DORk3a/zr3JSHclfUDbsoUXbc1QjHX6ub2lE+v3zaj9YkBSnbAc/35Vcjc
WBibLaFtRRAr0cqkGK1v3BQGXFIDVZXi+k37nXzsjb92bzD7XMSUSzNacZO5NbsP
pwFoR07XtYSZBlmBcwvKrUFzN8a4j5FKv5nNo3cqcDqHR9To2FUvnRpHshAf0ECT
IGLuXaTV5Hrd9nHxaUTJnS3i7abzD2b1ymaew9KGAC/y38/pJQ0ZxnWtaD9aOl6c
oId3lqkAoKimLFo8vJQ1r6M/wAWxVOVnXvhriTE7JiQWEwkl/8Edam2Qm9A04Scs
SeH9T1KsNAAHx0ePjqpOAJr1AWjUBJVMAZt5fgmKPXnIULc5J/KJnE5Tv3xmIENA
YmprBnzbJpGw0IlqT0rWRlqLX4cSHOQAnbffUUfRKub6lIQnvYGq7wrLFyZvBX3h
UmDmqsnQ9rkmvsHs+75MYFObc81Kxsv26KDd/ifFdwzUckHaelzDSzf/GMFKziBs
rVNBpTY4ZmhD42IRZKaxIXmIFG/VeEmeYDV4AN9ySWfFrfPBYOEg1I6gpEiaoyWs
5BKrgadjmijtHg3dcIWQ1iypykJkS8LXJdFCet+Z2HifLFGYkUfD/hwZEZbUxVBm
gq7QsLQiXZZOFonBgFzmzyPYMPBiBcFSgcDyqYbLaSr/1vy/IuvJ3apDgyB0jtbr
3ylw5MmSZTlM4srQ+VEeOfjp71/DXN0myMPPjeVMuNe34YuVnTP/A9ZLKs7DB2s+
54hIBap9yK+32I3MlyR/YTpVgH3CBFMdHXcnGTQtuNjfCyYU6JCDn3+/ZlR5EIqt
ZGENxqcsi10+8NroAjJSm6TxvCuN4dDlk47049oq3Gkla75Cyi8dvnnEr6Bv2EvR
NVwOskgimStdHLhhmS2koselD3XD04CZFZhlAAH8HsO1+1fMA6H1dOF21bv2XV5Q
CgCPuhFhabN2prDKQj6Qb7sXo9eKbrZqomP2B3j+RpdPF5AIHG4G3v5Si83r9RpM
HZxQVGYkEDqNRP/VAWxLe29KsJ3WihWrDiHoTUy39Ar4vEFxA9AcZ0wKy06RiFEi
Lo0FITCu+i2acYF3ugu/V9qy6OczU62ozsxy28CvXvDjRhda6JrA7jyiQ/imaRiM
lib0nZAx1AnSbiUPWAfGwOH6vr3hRcPK3PRsm4xoiK23PYkQEjz7+ynZtg1s5pDj
OQE5ruH9Fba3xINFriSkOcXrvSrAhBfp2Bhgq8sVLwYYIViV5W3W0nlQvBPnEVHZ
z7pXumLqhmriKlaRSGrSzy8kkldMXMp0HXiBZ8xyBv5ix3a0WUjNMNF8XcFA0BEl
YOfdMKAyzpT2s3xL2Qt1VMHA0C5IW7cwAC1gyCok3AHX4eUJQFWFSXCNP5VEE5NF
9jWtsjGZvfCUAEVvy24ARZbglym1O8NJCt/meDxZGMqaox+WkKSQcSkwwgVcuNUH
njkmOQFwyFMpqu1IX7il0esvn6wPZoMxq8RvFeoT8dGe8TrR8USyskUofChtCe1q
rFjumwVK7kBbynFCxb5KUzDpEAPzxkZu06hMmj+cc5yZAneMA4b7mq3itUuXhL/c
+/M+Pj6bcJm87t2j6SITLft1KiZ2bI5Q8PmPtCFAG/kcCK9yc74SxtcOWTIT4Q+u
iOz7wv8Nhp1FMb0KlbIfOH1Q14AUDD0LjyDnXLsOsE3jmyIkxmPRPPndxNndMgXI
CqhUV+vVHepJAlSwTAiDRTKRJATOicEmbb7w4A9EnY1v0dQR/wwPMuzirjCvGbfg
Tk13+ma7bIpYJets2PL0/EJ4gQdxsSeu2DkPYjvFzii5xd8sqrQRc8maOt5RLiKr
SSTrVp8uiF/9B2oXl0hvkCogX6KXUXLg3KyLK5craB/xHNyFBJXKpdSeC5aENr1b
cIMknvrcEqKmHPjjvREypcEiif0I7UCHoFZWsK3O4M/Ayo40WJ2rQnWirTIlfzvx
bTtIs48PpQnOAd+kb9A3HdlVVwDPBwW1fW5ov6PQNakNKSsiePIbGY/HTYcn1FHB
5I4Y2RcOxV2xXqPdQsM2OUzJFj2jqTNXFDf4GoppliE2GBuhiR95tZWrJ7B73tF3
cfPg+w2dvWlNX7khDFaNrLdx+vrWr2mnpgDEcqxqR2RHMlhpPwvSZAhMR9nZD/Ks
5uuDwSTtuJ0cG1FGYqIRzeZEWeaXoxwrSm/mVohWxyS+A3FL9bF29ExlJ+rWGwg7
hLRfwxB9hHU2IFLQ4YHScsL5/hyegw8DqU4tpNOiAVcK3VQdYqT1kkNHOmk+6jUP
2r1Xggxxq4RRCXyZGnXbxInxS5zx+gPxmX9ohghEw9684SUfmWvCbIRdE5adXBhO
s+HAse9MBuDnm9IcalWP78EBJVeZRiM8nPFJsQLnBSxx/WqU62u9Wlb0T31+Pq+K
kls24bIJPyT/vIcCmpuMYrcW364l6rSyyMu6j2ow/uTxrNiSlvpMeQzR/SRCPOvQ
fJ1fVjHmUzAKhHTGo15QaEqky+MwBTtMCYMFIGIHhqaUAzB/f15QPKJ91RT4dG9o
H+L9E0djYM1M4kHg0BbAHn5yilSPWiprcHsMulN0f8aQokKmgR+udyh0aG4teSMv
n49+2QkFJ8EddCkgo+mMuqXeN8EtKP5NPKJhejvsrxc6vJ0FEfUakpSmfqvKLeQP
/MKn4UnuGbIhITkvjs7fX85RAOn1VfRXQQCDNeNIby1YjyHKg5aaYKGslLSmlGES
4lxj3sk5poxp2krxpPygj1WDbtBR+1BOmuDJYKhtO8KWUTDHAmtq+LykB4RPiyzb
7thX8ymKFd3h5WFC0wDzshDY/TghQDtvMzIc/cmblt7oTmfuVwJgQZKc6zmVSTTv
yUhtL2iJQnvNWXXfrRxlhCkWPB0cfcNG61GekpnCLMJjIRIuJMURc4kmcRPFG6AI
rxyoMka/oajgAEkt+sfBzAkGUgLDnsyago3+9pypR1ID/94XKtGVbFk8/VPsovqv
EMfUU8Gmn77du7/bBlOD1rh8w/m8cYPg2D3Fc+mTdWK3seDn7oI5bSnV7LU3Fieo
/oVRhpx7JCcNBF/7pKQCFCXa20q7zIE/ESl1jor25NRB5kDNWLIRk+rrmLc/StIy
f+2LqAoqxwtj7Dn5RA2KP0MdomOySqkIOy200ltRRAlNkIs1C0Z1rUxAfCPY6x5S
ddscEmpFQh5TNNOzUY/E+TK41Ky9ilmQzKzwW0HEGVA0WQKSIMaG4bi9I/x/KXWt
ho3AdJlg0FPSwJYeohGKRQB1+IoGPBF5NSHNvpr93gNL4R4UoefFRDai6vuMbnAv
/AaBdkaW/dx9v2SrYDUiYOJFzLe5NIvfYP/554DDuWP8bvRvq2nMB6XQAGB1gvmd
zNBKLtXHxlZ8tfDjo9GDk2Uro6f9vIhKNa7WpuJ7ZlhGraV3uGLvomfUnmwqOGtD
EOyhcOY+Jh8jbTb9cZyrYoL629bfOpmTJ5ew/FdlH+WLUpBd78QN/qU3Orqu+WIy
HYLA9ZuaIN8cK3rEBXNtoWys+292si3Bl4H2K71gKCgB573vV6SFeWc3e+nfwR5x
txJpQcWIp677kQ+uiHPgrcO1YBINbEKol3tcFfUHChxx9kHWxb3SLurUmcRoV6Qk
4Y6dL/4sdB1VGWMeUYjjp5VrrcUXYBLV+jdbkkhoJ7/9nT85arAyMsDQAMpZZU0y
5WPL8yFDik94a9filwO8zbghCqFlWyc5BPZ6c2Zp/VMgl49+Co0Wv3CYzPlnU3oH
4pKWsBEHkm8A9RWlbsnH3n4HjSPRE71SLrQK344om5jBPISXA0ONdkZMG250v9gy
v+1QLEFA7YIRk4VKpntgUEPv9KkvYMOssHP4tydw8us97OMgcmesNdcmkPQUwBgc
RViOxy67EhuEv3lNjpKve2ivFaAlkf5K1FqM/MbnxUkuk5YVHbftDUFqg/teFJp0
dFwz0zg+jsY5kilRG48R6qjO5TmwmLVoko0RL1UOWsHugDPIOwCiMOqyHoJ4/UdS
FKXkw/gD9mZF/d5vA5NiihshVz9XNyK+jD6vwgN9cgUNjk3Krs7zbTaaVo8E+mug
GVqF+bM/rQpXKZVuFWlJpO4dxYk1ejJG5kMAOQuk2ZJotyclhp6jkwWUID+anWdL
58UwH68g+Xh3S8MKxlbbsV7yeKYSJa+JHDJkv5e3Jt1sK3tGsUCCM4dABl9OfqlZ
bIGQ0xWbwek3ddFob+s7nNj+Twgayf6xKAba3a64aWGHekBXe2hPv+ThWbmpzWe2
2t/mjeVyofmWX6XEbC/uZKJswxTveg9Vi5WqJZKsNCUOvxpY46vWnV/CKKQ0k98h
wN2KQ1Lyj+rF68BaOwKhto5xSENJCnD9r3bYGh7cuXYYKqXXeYb4v2Lb/l+igOcT
1cm126XLNIWBvM/7kB4LaubfeB0bPp9KbBGe79MbyQQo5sAJFqG7qDKQTLpYuR5n
uTn0KllHuKnDrdFTuOj6kXVFCEN3NKNayVyTckS0kHTQqIuA9bxz9p9LEgvTCmHy
qJgNP/9w/QbnfFGVZ9P6EFRYfWndQE/TOH7Ujk551i8L9W33PL6Ubu2s1lIR8ewi
4/+1TBb/RPFFljWfj4fBwhnrjH1acCmmAwwlMgYWdh7/dKzyCr3pppypAEHiTF/P
mqZwjBATr85XCOg6wvGsOoVVi3xxN8//Tyj6Almsr2UIHGRruTMKcDDWMOvKNGdQ
TGN70eWtcPU2WuRyBYWwmUK2i5cNS2KbQqoLfHExAta9Mg2NZNqvJF7V0ooVUcBG
EFAcKAfcZb7PjAFKrOVDoMT1gD2OSSVVUz56apPnVHTSxgp0y9tfAoB9XQ3+PYNg
+mCpSw0T0D+d+Qn4t0Ur2nmLyfe2ceJrBOsLrx5Iqxv//R+Clp0ERzOY+I8ZWuQH
NhFJxs8N5Vgzeg7UKfHR9LIrf4iDHqr1jo7BenMDhftjKwS8jDvO1GQyyskC+K0j
clyMGGuHh88Kuli+5hHSAMROqxuu6vKDIoFPKdA27/CJD9Fc+CiAcME9U7YvBs2f
6UjAykwDq0xhV4ycScbxPgFTabIoo9r9hJK6PwYGDSivGmKJVYG1WfKhyIaB92KU
wW4K7jU2Pqjoh/Q9MQF5MyDloCgAkOcG3RX34iqGznPiXzRJOd3ESNwtahPCDQl2
WlHwuqCZ6mlsSo0xNji/P9hVmqhWiWiReQSki0l0kwIh/nGvpW6rJNVQi7Nv9HdR
AoQp9mos7K/qcKYwrWmoAW6Y4SnEhf+E3tAVl0g1hSYgWrBjZKeG4emkLl0wgTW6
yFHR88lJrDsDDWmxNhKc+bpYxtinq1rO3SgZPQ9JwH32K3SeWnciFi6kZLDbKOLa
bq1TRf0Byo//HZlJiu+bzrNiFDytBxoz8YF9WxiDFrvvm8roUxEHT5TXgiN8gRHG
udsHxe93IOZjhOqQIzu94gmumv/9Mol418wG8brPCo+UAnxlan8Me1OgvpNRQSRz
BuT2oHxmGc83VU7eBj0iArgX2zNDCC2/7dCdwy31mhY/EccKXla78zlVEU99B5dI
TN1GGcTvYi8zQGkvRuake3QwBdfL5jU/B5WMpE2Jd2d93nGeubbZxNF+lDthiSLm
9KQcCWd0hY8WxR8Sz/3C9e1H/OT/d6eIYZAJXtH/VsQvorCkSOHeDw0ssFahQzu5
huyRRHekipfc70yU9qnxWkxFaJZuJ47zYrln5dhgk3JXeqaxaN21IrMLTbqVkq0/
j15Tk/Vn9bklrJVnwma+vBQa3lFuZgTEUingsoPyYasjKPa1qos0E+ZCj1NC35dl
xQ4iKaKpzxwr5xFaOC+RBl+7naEuRldj9A3+cPbNq4RNC4GGcgkoMSyX8j1wmTe4
UVrbpt/4aWQK1LHtti6Xa5tR2A3vjeartQZ7oLt+jxo6y8PKA+5bMpBy8wWXY8of
kUkcgPpHqoHxMFGsIXMz7TZrDGq9iezkdB2uUDrMhU6VJo8pwPtFvwVwnJ+m9owu
OoglkUh/V7JX+3dcdT5bGWCw0eKhDYUrr/zJY6ZclVKrPjfZVO2557rUGUV2fRMk
hWjVsBTA4oySR6+jlWTNB6L9Xc5EUJL88vUOGL1hpHlg8auDZVrwx0F+pznpUIgv
a6Jf4JBbwBiAOJ9dfzlXO6vxR0NMcfFRDrMeQgJO/gs4Y1zFabEMGCGJrwcAe7AL
CAYuN7LLN40KZiFMo8FQFw5B8oWZI4v5AZRle5nkGxtQog9w7e3AtM7la59QbEA5
pwgd7rQzSDNe9x8HlfXBE88jxoFZ2sr1oDL/PF+tK25MCA9Ic1RvZLgWUWs5ecJ7
owHHk4cxOlrGj5nRZiT0yeEN54StrGjNi1h99jLJBtM/HcMQaJ1uPxQ2JWdPhEC0
g1DJTU0HokMoMiKKdSImLMa91l1u1uUOXYeFxpJ7IHRcKlLW1HWtrD32Vd43CVps
hb/LZV7g6nsK4YT3Gy3q5OSDgBhn7HCIooqACsOT5vm6QSGT43dWrDzw6g26IqL/
1Z3wja5aIYM2SA9qcV+EL5figK4yFrBcsOBlMzs3bwJQxTu4qphtrsAMFcFij9gn
6N2hq1rkph7j9bvqNfosylDToqb9rBFXx5h7l22MWsrWzoIHUWEswcwNp0VUItcw
d2AbXFXXQLR52jAffkfb4jqbtcQ8OQioxEGSYKHeI5oMkEasE6/kThmDcIwA19S5
TkFNJMryCKuMNUR3D2ZNTbFutCJIh1SU/qsVCleNo3yXTepnxs0dlY8rAVVb3+dj
nbWwyQLXHe/sY+ZUgSPGp4elq1/OR4jWqnN3VAxXuQcr5aFTaD9X26EPUhgJIv+Z
LvMLHL8ARpwh2FV82Yeo2SaLryj5SZNKlk3UZ38JTr5QRI1WgkRHrrsdb++6y1oE
ph2s0rBPAwgMihk3JRKyX92iB7sFmFRf3o44o39kC4zqA+RL1wMnr0WpvwbY52fU
alWbipiTDbXrdCaRaGKyoVb/sLskB+bf2FjDhoZJ2TUVdVvW/okcxgIVbZWfWNlE
Tn9UIRJGJgiIz4tWgK+dWXJB/yEjlHINP1+jS6exyNUhuqBp4JDwpMxIj2iC/6Oh
vLNM9oYHiIGV7iyzLn2a7sUkD3wIqPlke+H7+ZJPUZcVPBjTyIT5FNjItfBU/ASW
O9QOWjnVywkdS4wq55vt1mr6fTBaBfZ8qkiz8a7YhMdvzv5QKnJOAb2SsWsVOKwV
ko2W0AOl5jcjblmrlUMe0STRp+ZBo3WYjpCSxukvVatXKk6dC0A6aiBkdMLvZhsG
w2y5Fi/JCkNwlGi6Ntlc57332t4fGN59XIXr5grwcivUpSRh1zR4bJB6ffXas9pA
A6T3loygIigqrg//ULwLtlenu8OcNJUgbFgcFpMa1nPN6Bqs63ozosC/Vs4ksBI+
Uk4SsSe/qiuhokY877YvHk57Hw2XQ9Yn60Xa1G1hk542YsMoLC46AMwqwNzu+0Yr
sQJ1jLXpBfIsAy2sLCEzOTYbSNbQ9tcUfW/4RfjPVdxTvPu6pxG9kXOvkT9yh6J3
nF0j5AB77j/ihKkGG0XdxOxIJuGhNietkxtfGVWe+Ovvalfp0g4k10yVMjcw6BlV
k6ZX45N3ZG0n4LiUU+LZFV5WQ34SL6ayW4qOyOgWuR+f/diNJODdApdN1G3vvLaf
7n5u3EDDa/XLLLIPEPowfICRe/Jj8UhwbCtgVO4tPJUAKsin/ltJ9/hbsuJ3Hta4
FZjmibPyqguy6rHZH86O7ZPrNelajMV7zuxkeBtjIlerjpje6k4HPWhd+XCrvcEq
fbPHFeqxax0dfqKopeI2/kugrm3iOn1EVfZ56hiGmE8F1tcl8DyzuDwA73KruRcU
SIdCJv0Aq+4aUAJ7K/no3Bv7d5IO7kuJrprDauWqzkhC2kp5M+mZtskQk2K+h0Ro
zBRapSr9bESNGh1glh/nUuNtDxGXoU06fAFqLEXUEIIQBqqhr40GYWpq59ZkjdkR
qf1OI7iuP6E5OTBr8//JCmmtau+jAKMlNzg4l6AtnD/J8PcRMVDF+ottXz+yJNXe
zm8P6Vgz3quI7CtzRUbXbge80kfX9wHSLDffZzy65pgP4i4lY/CJ9xmZxehxNfmn
C5Sbq5lnlJazKKSWtVEZK/Kuc71kEsVaQajQPdBT9CGvkUZCePh4UOVAu75Uuz2m
0j7Uyi3XHCuKj7GTLxC1VG8bjQujcTeVkmE7vQlWnoh/V+bOkMOnrLBeC5Ki3rXC
1FbZ8u5hG7fUDA6rvkgcFQF+/atfPvZyseSDvMEd5fsyOBt7pyxSfwLDAfn0lgcD
WClKAYuj/amHVtH5/n7g1KVYapej9dJ5yhgYxFSi/YnzXczccezkeyINMZ8eseHH
JbdN0uswx6JOyvmSE7VPxWbYk4PpN/AGTfZGmbOYrxWe/tz0uHefKGwSGJcyHUGL
1CmOtmH1T2VHFwOUZj/PEc8Llt/EaTrN3d+N08cWeHm/j9cv/kKwxoPzriQucz7e
8QVQGRRxpqCdzq9o3G5tWIYVsc2GTK8YloupZxdcrmEvOgTGb3TeAwcQ4/p7jL5O
tiEvVP9ExMbf0onmeTxU+CbkhFXpmvf0YjraGg9h8JtfCRuFT0xWaXX5imO/3CMW
Z7lZYDnguWezxpoVGaNGuceuI9hqBJNKeB7HT0FK3usO6zkllaHVkcI2+h24qHuY
ODhbWuom3PlS2OONcdxv6hVbD2qqIRM+dkPuWQXzCw1XwgNwplyN93QybUrSeT0c
XW9FPxfijPq5wy/V57/7i5kd/BxLVuIDPu5QsXMP+KIbNrb93aPyekFUQiksuuvM
qjlZTKUnF/QRhOuWInrlfmjy+q8bK42uCySbajqHMbYLDiI8LJW5SwAUxlExECaY
eFOiftzJny8OWS8CXbFbL3BRyAvdYDGtQ1OX/3dwzm3V17yi75g/qpu+ulbJU5Y1
ApvhWp2gdSbuQiv5XrEcBqHgo4R5yMLWFUgStPLqB0+E+kNJxFVDlkov2kVOT4a2
JPfhUtNfTj1DlN4BmMWPBeuapxiG/dQHAAQNDmzF2No+J4v2tuhGtTxov3MAEEHi
MTg7wOPBfno24rEFPa6fFS91FBdyEeFTu4OSjHTy7Q4hwWKygiWK7zGoNx8OXH6+
04MvsGVPYns/CzzSIqWQGM+5YGjtGwitMYLQquC0vjCTpjzexPc0LXRrNFPYeQv2
EyYW4oQ3wvg7O0oSbcHbhhu232zklTYL2UejuKaTNVgGqJa+yHpGNGfVk8NzjukI
NKFBWBAB/0mRuF+wJVVCP6WEFA5hW/e65Q5x9YsD5qrBetFIJZWDipY/+zAoZtSo
C5Wqs2jEVwiExACmhh+itDHMAYuXdPSMhKY8xDXw3GkL7NN3uXmGrxmX5mkkVZ2U
EaMlimgddx26MQtRIL7i1EFnSmLaev/1u9JE3Fjb195lMqMHoAeApDWnqmMCGmkY
MdzUz1dX3XZjLbdpf0KSm3SloRfoqqd/J+xgNK+pAn7kXGpgPdWsm7s4nRd9N4wo
HK/8If4i2MMnBWjb0FgkGZA4i20WSfaqnLmxHhzukMHvsiZUZa/DvE7iiyLS31dX
44z3mteESvRQEIBOJN+tmZ6kz7MpoLF3hcBvOoUCd225zernHyl6IFckjrhqxArc
jIB402xxZc7Ig1CHpT/+Jg/9xfsL42gnpygin2BackTz5phTbrI2XKVm+mfCiehw
CB7UHhszc2sCCU+xwrGzNuWlYRtnW5Mci7WPg4VKFHINuH2N/hrmsvjSIRPyP73v
cfMfCzLB3G9uXmew97nZUb4UKGiWcMJ+LoJiZENfK1HH0Vctfa+0oojND59ReUkh
UjlNGqnW5kHGnvOQ7ZPus8n7M8qNXEJ5mv1wTapFjvbUr0vtbqf2l4iJ1qel0NIr
kp5zehNyVNuBhjg8U+GUI6gomkLkPAB7oCKBELvsuiYwB8WY+effjnO2a4cuJAL4
UOJDIO4DcsNOVSZm5nPsF35v68U49cQkGFxPx5r1vqNZl5xMNgkP9qBU/djHdZFh
epQ4/mCQjbzBtT3/3c7BGQ9E6lB5/1cNW0OnpSVUIabgq0qJsrLeMa5zfFR4djuu
6HiZiM7xh50I+dEm+bg8Trut1TfNc6KERGPPFL1fZyrP+7VvoGHr33ln7+78srwl
YWKYKTje+DBqtb84pXCc/7h33oYMox55QMjO6r6PFGQBIjowOAWXkTF9P7pi624T
8VHMYL4KnkMs9Vm0d+ErHHZsh2ij9IX2vGEHp5baC96WLSKYVocuB5OMcXLvAVG5
clAn+G4ufaweffne/jVJ4ubd3qoMIdx62DMicMZ5OlWW1CNfey/zeD6xDnvnxtIG
uwJVpl6wql2c9LKPOS42o8rBJCUYU9z2RB7OAkBZ/T3fWIivaSYaFrH/aHXbyjiX
hU4Qmlepr34HviL7IT3xPh3ZQm1iDTIgWjbL5fqEF60Av/oNodNvfH1EyMVPMWpV
lQFUPQd0A/05oPZKKNVRtVCjva525F4fRPNZ0oRlDHq8va5Wj6vT/Gg0rd5Qr+3m
yn9F7QOTgBVFVOnrAxLQg4Ce2IYTNRjo17WH1Ctc+YhfqQEtfr4IV3cHZyv5jbJA
N3445g7BeQKw6L2t/N/SVzxS0HAMAozgwbhWvHZPEBDXtJ0ECXdFo9i+aWaqL3cV
30GeRIh8JSw4d+vu84fTYMNf0lDQ4ettRTriq9ZsqilfjBOULsbLu8zE0sKA2aew
qxzIP4smS6n8s6BUJbuazgEtE7i3U5aMKn4FIIXw8PJ7ceY5gtYn3roQiptZnfaE
TQ39mQNbraXGLMh+7uPbsDQrlb3YL8l/md3SdJCsH4v/yJhec6fWAmKuSOyAdJmZ
D1c+ncHzACvCA/pYeIkxirKVK543AimafwkaDx8ItmlBnKqOOeDx/Qcs740o6Hbv
hfJSP00X/GlO3PumuzjFqOMw6gtGMs36Gky1vJJa8oHbdUTOgz6SuffkSaMeldF/
vHX5rLdIzB7lU4wqdaDOg6DlJnm/esbf1jaMfwmnKqXV5xvP0jQtEAoMhgzN1hLL
HJntn8m4phySfyMiwvVsTqGf1JQ0oeeb+rVSP7KBIU4cfREW1RA15ZqArY908+8U
Cad9YCdEkH/vJ2cKXhBPHLxOb7EnFKKGCBZL2o1QmBxB4qXEtg3Wikcd7IrpG0HF
iux86IsYgPX0KwwzC5+lNz2WY16ZMOJS31ccGFPz8ngToUeFPxGsD+NoDutmHQnV
rjhbQyZUN0fYOwMQFyPsrIKbMEA2mc7g7/4Z4BkM+wR+T2V/YEBJ61jQxZtvjRO0
DCBdHeQVYRvX53GcRgT6T8L+Fg0hQQOiL3s8q4eNlWbKPbG0+5juVU9fkU+8kyEp
sHQcZZ26DUeGi2I/trgcUPjPQgmyt9PhN0lHiSv9nOqVZTuQoFBBvaWMLVvv2Qb/
JFeBRgzMa1/95eq8lwzgVPgGcXOx1w7FZO8k3/mVtxOziCvXy2knYFWTtIJ0TPno
oanh0LxAmuq0o9V0UfIbqe1MsYmHu9tWg9YncminHcbSI8ptADs9xkOhfEiaj+LB
jJuDid47u31+K2gTdoZRINRhW9AkOVI4L54CGyzmNafXGOJZFYumqhHXoduc81iK
McAX1kNtaEUYbfjtmojFxZEqAK7pBW4hn6ee9aV+51Dv+naziskM8RMjE2+9Mk9R
A/uW4xy9HXWizCyt9wMqoxd0nDAnCRs+q8/La7ZiZsc3HaPrCMkhvGNyoBHevL8E
z5pqBvEcqbUG9YI6522fOtThcvRvoOCjUJOdzqlLdupdu9PCPVNHmcKKNmwtS67Q
8d1gHJw+N7zgPnKC22Cf+9QQ88Y7lLUKqlufwBfX/svor0f9STuv+jmSGcUQUGqh
mqLd7omfUDJNiLj6p/EOr9Bs77oU3wfjPlYJdOGFBE8I/ZblNZsBTvf63sQhMr2f
rWQe8IDEOFRogACE/9+JE+gRzgFMaOsujHfNotxjud6pFor7p2XOdsFBvofqfk5p
bTGGP5wmGR/Ji22zeMCy3vDw7ByShzbomncbSUuUajM1QOoq7/KRAx8v6i3VmtDp
HMOpLkFKfa9j520GBaJ7ELh1JdmTAd03v1Dzx750j97pm89Q/za3qXoLDocT7g/l
mHHE7UZefdnd9k0+wzoDQkgGsQ24+fLtNVG5ycbcENkmXIufB/uTg0h3Vd0ZKsci
80NSTl1FM86IMe2Ez5I0B31if5Xom/OyaOxBZfGgnhzsOe+NI4MGzWC9nImMuMI9
qPa4m/OCH3TqVoKR72UY4m3huzVEMwGvAyZXvdG4ABhnJar8119hq4CQwURKAlzF
estPkrji5TSkxSigcjUJfAgvJrRyeF5ijessY68Gw/OHmcPZPXVQSGTIe9Ghp9tJ
IaKtGk+ZRZLqgQ5mZrGO/5IqclAub05X+JrOo/WC1swPbqCTo8PIF/U/6yblKIgO
eDapEB3+fBcgz8Wc1ZnOBBhJn93qZ0gwkuxmgODCtHSMOIJFYInL/TsVTKQ/mMiL
t5T15CFLWuXvIZm8XBjqo2mTrUbhnVQ1hvnb32LDRk9MXXi3N56K3LAJ3T0JgYmz
KaQoGvXDBKxM9rKF6L4D157AZDmzwMv6Bgzg2crRwIiDhFA4TyYOUnoyHPR8SN6e
QGrv1bvs4bVYaKoiEVd6xqHKlThYIHGPh6AQSejfdwOPfErJKBHbaw533diwMVS/
obiobmOpdOvfSdzbdlmaVB68JyTbRtF8TwH7McZG3Z0bTxmJdL1FvP+0EV7RZeWS
GHG8tsBNdnsVVNz3ZKoHTmoIZpaAtJDCam+dTpvFhmeDbIQr2rf80kBK5F0QvMeR
mNxCUJ7/l5uf6+vYlh1twC5JLFnZ8u4tCGhcfoSiSoBRMHoLnYFGwDIpQelbbRSo
qfOiSdVI8mHeTPbuzbPqRWri2bSCd/VVAoxkuvuJM94xp2Fh5J1RC8u5xZXuezAU
UfItjJOV2b7DMl4mS18uW7A2rkGzQrDMQ3SgazAArXdZbGJHk0e7YiI44h7v9X0i
W1ALiaStzZRnQjNIuPfIQqRsV9l1lF5Vt+kB7hK4Orw18lGyOmuiwory+59c4nqI
d1cGBfqg1mOH5s0kfZDNNm19YDmxPDSW5Xs3hV7sEU2d6ndqenmHE3eU9RCgfD1E
FwZra85jixwXK5Ue4oXGo4PfViu4eQVLXo2H4Is2neTzhbGsD/+YCNRzvPjCl3ak
TTQFk02eFqkFgEr/LGQnU6fywzlvIcelYN9flnFqcUN70m5OHHuX8GxSTd8zpTKk
fdTn0aYxmWBUQpI+xWFFxs1NOir8Ok4Oea/MoMLBcgN8Va7KSJuifyX8crI/oGLQ
eXbJTiQeneGY0x8IeOSthKXZPIEJjww+YUOGv48OfxtjnxfOosvp1L/FpVtNLkHt
8Q89jpBnzY1//Rlw9V0NrXt9kXN5ca7PZZgJREROiobbh4yuM5FfEWYuLsNtPSeh
ujruaK+VRp4AovblQkmHEN5hxpBRjn3EDFMNCtxrPnYZXl5nYo2ndeB6bCmDXRt4
fHY/ye2lfCrgct3klvRmT5dX9XBy3Ku24cdWNnvqZIg9c29sJDaT5ank0QLoTibK
ybcL5M5TsfPrGyN0LL9HUJabp+EzVmzWJ0g9onxJ2UcBUoGy2D6k/qZWtBfdPzKW
SG2luRF0Bdb1xv8aWa6mJ0QaI5hHLcxZDDawEaebY2OFiUHxnofKffBOxqsF1QXZ
oEUIR2kJr4V3fROm8hyGQlkFW+0ToJsQr8kb6FNigrwlcaRQAWUvcxiNaYK3Z5eH
Ptf5/JKBzK2/9YZJsagwJ1CB6+Fze4DdilCa42JJJSQf3Gsrol/adfgbpLJVm2X4
HtaK4rLgHJbbHudedFx1iItHyHTbPtKarh3psj+XHjYzQSUSzrzvfzRG71G7x0Ia
2LgdxZ5tBn9wDfCWOXPIklCFz3Hc92WiG9wbveIYS9oB47pjaK8ec/1H8JmP/AQH
xaDswh2jtYofyy5/ito9wV1JNFnWQRue6xGKH6/kbK724o1+xmpnVOWOwYPo2Hwa
gNpQ18vk/kuwH+R69umyUm6pVnKykgytJImpHF25OnxucPmOVLdB8H2pt/ifw0rM
3sY9Vxp+Y2eHDQrzWB4+gYcAl6AIrpteL2xIXmfHfHatXIQZpjjn7U3Y14I7+ii2
OiLMUT1K5y5YhDqoKJSuAEDHSJF4n5C92/nyFuUF15GEkF+bCLukrNZx9+Z0iZrc
kqCusFEG+m+HITDcGPEf2PeFE9wBcL/E9U9pUiEdaDOc0eSOJtQ9LOtLK2M/Y6pi
E4eSlOB3x2YLxxLXqAYcZiTKnxcyOCxwF90iFs52kd2RqEkqAJYOVm0p4xlTnRCs
2GIMsfCpTivx9FAYI8qmVhrpgwIazCgwv3S0yZRdmZ4vhSv7u+1V7RpB2AOq9w3Z
67tAP823XktT/EIt0JkMUQ201mk8DQ6N1pOZsM4cJ0PIquOxSULyeKvQl/avvFA2
lA336+IcJrIsMnKTiraY/wr+J4JzVov5aUyzMiko+J3Cb0E6yyFqzS5ghuJJa+tr
O+UDgD9IbXpcxRqpjn5dVopF2i6iYwj4pLQNJMaoQYkObBYi/KeDmxsro618NhWb
rGoVisBXF5F0r0WqC3n6b8L/Ta9ZMKhMwhDfRpVcxjNyDTcAjMinYjIfw6WHB35d
vaEX9vZyRfAUn7CpEvFDZTUx5FZ2tfIgqv07b3kcoLSVFjyHQylcCOijv5BINcoq
Rxpl9sEPksfvKi3yoXmhQLT6F/Ihx5FyHhOUIN0uHAxWeofVGMkcpZvZMmlGE0iX
6iTMJi3AlKFzvpucr54fzHbT9GCavwdcSmsS9uQyUyQw4zOsNv1qnPYboy4JoAbJ
33X6/4TUMOvtRaq/+lw6t0DtD8rWKN1fG2UJ/0DGH2PjoiNqn1pD6ihKr6c2JmTH
e1OryJN+gdw/7vX40PPWKJ99EdayUESHWVGaaMTGUjw41GmiryzQfOT3H3BQvq72
Xp+2PL/J/HUIRLBlIQFP7+Z/HeR6BIAxCcIXdSCfv09Ud1F+tg3KNGBihZBMCry6
tPfVD4ZQC0X9JwcWCeFf98I1UfbW9nLg1l72bH/u+Abgd8Zv8NK1r0Qx7FnkRtqb
lj/bWK94jrrzcVBCKpno/RoPblZPoowvbRTWw9zJ/kG+cG/2J4O/tO0EKjHaJruX
XN3TseZXbf1gpjlYvTHkKV3uT594/qM0g31B0wT5kRlmUTH978WuCfi4JokTsKMu
8+d0qQBFkHdiPRaC9l345AwdSu8sD0XXTqUOgvQc1AEkMOC2v3xbGnzXDV2ztvaY
2seW7VGjEvGfVcgYm7WwoxtujTM5/0TC3rFddOsBwpiwNwMIn88S3Xez75b20BNr
+3nQ0b32Ky0RpKoEw/fkA7VVII7HxSSM6i29MlhFDs74iwpTWPT644Rqdcu3xT3T
oRqdyXfM8jxGi6/DPWT9ao7ks7RNQultz/OPPTVsA3YDvcOYnoi8TYmUrqvyA+Os
0UHC9bYb+co2LMdjigeyFLWAb1qtuD6Uut0n+mjHRHLWRe4WSpVkA4XKsp5I4NVt
5zuGvpP+SnHRtCM1I5gP1C897r8gwT2ZRKskA2amcWXukAMsZPcdkng9mB+8Zofb
Ct9ENccJ3/L7Kzr/qfsUXh/Yshao0cTUVrvEaaWwsaSSdDMQyIfC9YzXxfGjgaxm
eWucdshYzvI7IL67ARJ47CA6mW9niTJ0qCShTjqMFKJeqJ5BA6yvr+etXAdh75jH
HMyxMe37XXfO7Ee8z+xWIr2U9U7qY95ASzFJXJd8ZfivcJDFA36Uf3+XLPBJpfqG
qsPRy0W6H4MHKcQSuoSomaQ05ijtI1J3pBbyKcO2luW3tE1lvBWhq6pnUeRFth5I
4xhaRCeoHP81lQ8r4aARwaq8tQtnLUn8ojN0WQxx8x5VBGYaXtHbtdpWNF0w5M1h
rJeuh7KGEu0AjA6FKllzSOwPg0vmI5QEZpE+G5q6nfi3fu3bcAX6lhMCy3ko51av
+RwUzHJ+S8UaV8Dq53TZoHk3brwUu6Vr7HXmWKy0Yi3UHlHIK8cfnQNYqcjvjUs6
KQ/asp6FWtC7VOu8DOnnae4WkyU1jvNjeZN7+y5OYj0ME7rEVoFL4mAjQ+jFDDdd
z2wHiFpa0jX20YGZMU7PKQHDlj0zzdT5LROXVm5vmI/gqxPG9LH0dSVDBb6IQfUD
EuHDoGuBeWb8UBRfl5FH58nFqxX3Q+PcWHaLH1iMoNnSru6o3iKIr2JnVb/7CQ0k
WGCBNbuBfIANDXRUPfaXxZQ+2/lMxsquC9fB0VS5OPkKd5FCqOCUi5EXtoEplIR7
qUzcOBq+BwhiWiYTbssm14ipJRHmb6ZQw+A/ZRDbCbioj7gubKAoWrphe0b54S83
re6c4so2b5obNWzzg0LdYzRsfZEXFuymIzTaMKoW2v0I0gSZhZ8J+KJvjHWo9Pqr
G8wwMvAQjlVIuxELP7oxdh7xnQ7y83WkibXBiPz4KTDlE/t5tUlWaMoqyGcytSFA
sTy5O+d9EohzfxVPgcHhx647lHKaKOJqHWbGhxsPK555jVTWGfYcWl5r7uphlBlz
8kd4gAx/eO8yQxkOEO25linXUKYik/zBU6UQU9n4p1MCBI+oBC/RT8A2B+ItxLQL
rZiPYjFeB7M8jrkx7/Durx3Ix13oBV1nOQFGV2EROhUMUK0/NFkHi+OACth0JnPk
gnuvgGcMoAKo2QkOvhojDc/zn/Eo1pSMlEycyDSkoLF6xojCI8wnLDFxHIeMWNvd
O6VPj6JlbKLnstOWxHzz8w66octTPVWR/ZgrIWZLjMO2RAzG0Wjw2bXvdE1QI4K/
aAKQnDdURU1C6jr1eqijW2+1WleIQgE8DCgrbvto+L79qcaYXuyE4aV1WDCBYpAV
Wy1r4VilBBEToseAK5BQ9cJOqbAAZUesusPORGqGNDLxPX+8L+6KlkzNgjYDXwQG
IlERKhBmjeKW4WKhJv3Uesuae0QlSF1ypbnwYAnzAJGvJe5bMdzcV2obdB54K8SY
6rCJ0494MMnLusFa3GnKA5aoMJemx/NdhOV4Le7LNRnbWE02vv9uKDguSUi/bnNs
T1g4FbuuVtK1tX0DAsfRuEUbBDpKHyWhh12zUN4uTeyQ2abdEWhDur80gbi4rPTR
dd7TAFn1kf/Aq8amfn97Ul3Qv+hAm9C04SmgoDg2g2Vhs/byanEMVR7g+QaXzxTU
uuSS4VwceVt4qhwTSFLrXaYtEIWCUe28EyBG8l274yqWRJZUjaUnMLku9VhJvUAo
f1rL5abH9TrMwvrk+6v/vX4mwSCjdW3RXY4WAi1UrXsSXRupIRZtH7o1RYGaUiEy
fWCQUNlt+w1SAsS1ijPdQL5mS3iPGVKtybh2MmUnK5wgtopj6Ku1Pqwaoo27GxOd
8mmAZrMCzzJncz5BlntqVMoRKSp57G3as7BOsWule+epacvozeueYR5uByb8kzF4
h+GKnWvkLe51UODQprwcUZPSdbMLOazgpGEQJJmZPkEQsgIG6kOP0TyD3JIxVpJ2
S65yUDgbvpBs2aZAF4h+tGYe3DI24WU79F8qAXb/WEtky70/pFFRJRoL7v6Jeygr
BD6+UWRqU7l8ozDRy3cFNmJiY20V9GwrN3S+BCzr6QLd35Pwh4kbn2CdUtPedEjW
ow5hhndMxoHzqLsuDPLI7TgXUKKsAUQTN/sXeCE6sOKshh1VTUotbjK20pdFT3EN
+kxfKMgtAEuWIMEPgVJzGVl44mTxjb7f6aH8F17beNdEH42uNG3G0v/gGpbeY8Qh
qu/uLfwPs8ZJ1Zh3ewV+tc/bPK3SPkYY5XEookN1Ua1VfzD3UTy+EgpCRu/xXASD
pJmMC3LbE+Zd7cEctLyjl0fMDuiuYfIn8PP+55L9eNakGqy08xQl1mLuuPf5UCkg
VPmq24+KHDdJb+XYXn/oKxiOxLSDHjhQ5u9PBzTlwhHd3W45frO2PLB72nOBiEc8
iOPWGz3FtyMOZ2sCysPQoH1QAfubHtQd4XqjsKQRgdnh27aSUtPrlnoGFD80zBOc
s5zgEg9JiRhgSsFmmuq1RGH22TFFns+4rcmV/odA1jesyBQzmO0En4TUudlllacE
G8T5vTdtr1Xbghpeh/VcDtFrAAvTLQ5DF7Ibm8yGUisHFytleGaupDhXmFcjXw66
Z1KJDQ/+EPSNNT+Wo08IdIzpfb5q5WcwOYMtJnx5WTd3H9BlPcjo56bh0vEzn9mG
P1+T2gzl8yU/5EN8n09Dhr5hHIQJabuUpE1R+a0lYI+vnqHlOsV1+nQdPlZV1M2S
q4y0hWoc9LOr156I2faUWFbtpKdS36AlGgIDSRLmn03Uvhj7Jw/A0NY6rhcwR+Nl
A6XUlIapMXOAVNDbnnIzE6jaH0ml0vLzyIfUzwUnMxWElRMtKSOWzcehhwHK2BwU
jG7HQOjnZV40LPzQZ5NdAShXnS+2crZvAewtjVmzGhHyKo2xyDSSBpTbwepDmJRF
DtCi8Fo7zbeqtWQLajvppWJfEz28ohNO9ZpSHhOCuQQCI5gLI2TpGpgJohstpUKJ
1Z6O7HVaIg4ERkK/yZ7dHxCL5Tk3Vy3Sm+G4w/U+WtoePlm+fI5prhR90LzB0LSS
6RcTN7TnkkBVv0iFYjZutT1BbA1cvlAd6TpeGN528J0EUfQpov2aSsXZ/sjyxElF
2MUTmSdiTwKMx9toDyYLmPsAOUalvw+UxE8SRphAMR+LHPUfAHoIvFI0FMhrxaQq
7TV6eWXNfDh0ONZBTfy70GnCify+9z/qCclfQ7VanVexaKiJFoWpePrjGeDN5+cO
ENAwtOXfJgk6VRrGWccOqL/q1D9V6u6OTRnl5ixJ8ZO6rCfGVDqcp6lp8q30JWcr
Qf9yPkjxa9cH5vQ8MzRWmY6mL2C9yJ9w96le3y25wfhwYfeagdKbCP7faMKn/Pgq
58bCLBPDSDrV08M1jkv77A2NNudfje82nE1yHQMjBvzjwVa+we8+foKXdI/jkB1Y
5NjpeKNXLwrTxM8+01/mFdz75VTi4xAETXO4MZZLkGy2VlX94O/sgRaUa7ruMn/x
`pragma protect end_protected
